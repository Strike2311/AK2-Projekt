module PPA_adder_tb;

	reg [5:0] a;
	reg [5:0] b;
	wire [5:0] w;
	wire ov;
	reg c;


	PPA_adder adder (a, b, c, w, ov);


	initial begin
	
		$dumpfile("wynik.vcd");
		$dumpvars(0,PPA_adder_tb);

	a = 6'b000000; b = 6'b000000; c = 1'b0;	#10;
	a = 6'b000001; b = 6'b100000; c = 1'b0;	#10;
	a = 6'b000000; b = 6'b000000; c = 1'b1;	#10;
	a = 6'b000001; b = 6'b100000; c = 1'b1;	#10;
	a = 6'b111111; b = 6'b000000; c = 1'b0;	#10;
	a = 6'b111111; b = 6'b000000; c = 1'b1;	#10;
	a = 6'b111111; b = 6'b111111; c = 1'b0;	#10;
	a = 6'b111111; b = 6'b111111; c = 1'b1;	#10;
	a = 6'b010101; b = 6'b101010; c = 1'b0;	#10;
	a = 6'b010101; b = 6'b101010; c = 1'b1;	#10;
	a = 6'b110100; b = 6'b000111; c = 1'b0;	#10;
	a = 6'b110100; b = 6'b000111; c = 1'b1;	#10;

	a = 6'b000001; b = 6'b111111; c = 1'b0;	#10;
	a = 6'b000011; b = 6'b111111; c = 1'b0;	#10;	
	a = 6'b000111; b = 6'b111111; c = 1'b0;	#10;
	a = 6'b001111; b = 6'b111111; c = 1'b0;	#10;
	a = 6'b011111; b = 6'b111111; c = 1'b0;	#10;	
	a = 6'b111110; b = 6'b111111; c = 1'b0;	#10;
	a = 6'b111100; b = 6'b111111; c = 1'b0;	#10;
	a = 6'b111000; b = 6'b111111; c = 1'b0;	#10;
	a = 6'b110000; b = 6'b111111; c = 1'b0;	#10;
	a = 6'b100000; b = 6'b111111; c = 1'b0;	#10;
    a = 6'b000001; b = 6'b111111; c = 1'b1;	#10;
	a = 6'b000011; b = 6'b111111; c = 1'b1;	#10;	
	a = 6'b000111; b = 6'b111111; c = 1'b1;	#10;
	a = 6'b001111; b = 6'b111111; c = 1'b1;	#10;
	a = 6'b011111; b = 6'b111111; c = 1'b1;	#10;	
	a = 6'b111110; b = 6'b111111; c = 1'b1;	#10;
	a = 6'b111100; b = 6'b111111; c = 1'b1;	#10;
	a = 6'b111000; b = 6'b111111; c = 1'b1;	#10;
	a = 6'b110000; b = 6'b111111; c = 1'b1;	#10;
	a = 6'b100000; b = 6'b111111; c = 1'b1;	#10;

	

	$finish;
	end

	initial
		$monitor("At time %2t, param1 = %b, param2 = %b, c0 = %b Outputs result = %b, c6 = %b",$time, a,b,c,w,ov);
endmodule
