VERSION 5.3 ;
   NAMESCASESENSITIVE ON ;
   NOWIREEXTENSIONATPIN ON ;
   DIVIDERCHAR "/" ;
   BUSBITCHARS "[]" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

MACRO PPA_adder
   CLASS BLOCK ;
   FOREIGN PPA_adder ;
   ORIGIN 1.9000 4.0000 ;
   SIZE 106.2000 BY 88.3000 ;
   PIN vdd
      PORT
         LAYER M1 ;
	    RECT 0.4000 80.4000 102.0000 81.6000 ;
	    RECT 4.4000 71.8000 5.2000 80.4000 ;
	    RECT 6.0000 75.8000 6.8000 80.4000 ;
	    RECT 9.2000 72.2000 10.0000 80.4000 ;
	    RECT 12.4000 71.8000 13.2000 80.4000 ;
	    RECT 17.2000 75.8000 18.0000 80.4000 ;
	    RECT 20.4000 72.2000 21.2000 80.4000 ;
	    RECT 26.8000 71.8000 27.6000 80.4000 ;
	    RECT 36.4000 71.8000 37.2000 80.4000 ;
	    RECT 39.6000 73.0000 40.4000 80.4000 ;
	    RECT 44.4000 73.0000 45.2000 80.4000 ;
	    RECT 50.8000 71.8000 51.6000 80.4000 ;
	    RECT 54.0000 72.2000 54.8000 80.4000 ;
	    RECT 57.2000 75.8000 58.0000 80.4000 ;
	    RECT 58.8000 71.8000 59.6000 80.4000 ;
	    RECT 63.6000 75.8000 64.4000 80.4000 ;
	    RECT 66.8000 75.8000 67.6000 80.4000 ;
	    RECT 70.0000 75.8000 70.8000 80.4000 ;
	    RECT 79.6000 71.8000 80.4000 80.4000 ;
	    RECT 82.8000 72.2000 83.6000 80.4000 ;
	    RECT 86.0000 75.8000 86.8000 80.4000 ;
	    RECT 87.6000 71.8000 88.4000 80.4000 ;
	    RECT 94.0000 72.2000 94.8000 80.4000 ;
	    RECT 97.2000 75.8000 98.0000 80.4000 ;
	    RECT 1.2000 41.6000 2.0000 46.2000 ;
	    RECT 6.0000 41.6000 6.8000 46.2000 ;
	    RECT 7.6000 41.6000 8.4000 46.2000 ;
	    RECT 10.8000 41.6000 11.6000 46.2000 ;
	    RECT 12.4000 41.6000 13.2000 46.2000 ;
	    RECT 15.6000 41.6000 16.4000 46.2000 ;
	    RECT 17.2000 41.6000 18.0000 46.2000 ;
	    RECT 20.4000 41.6000 21.2000 46.2000 ;
	    RECT 22.0000 41.6000 22.8000 46.2000 ;
	    RECT 25.2000 41.6000 26.0000 49.8000 ;
	    RECT 33.2000 41.6000 34.0000 46.2000 ;
	    RECT 36.4000 41.6000 37.2000 46.2000 ;
	    RECT 38.0000 41.6000 38.8000 46.2000 ;
	    RECT 41.2000 41.6000 42.0000 46.2000 ;
	    RECT 44.4000 41.6000 45.2000 46.2000 ;
	    RECT 46.0000 41.6000 46.8000 46.2000 ;
	    RECT 49.2000 41.6000 50.0000 46.2000 ;
	    RECT 52.4000 41.6000 53.2000 46.2000 ;
	    RECT 54.0000 41.6000 54.8000 46.2000 ;
	    RECT 57.2000 41.6000 58.0000 46.2000 ;
	    RECT 60.4000 41.6000 61.2000 46.2000 ;
	    RECT 65.2000 41.6000 66.0000 50.2000 ;
	    RECT 70.0000 41.6000 70.8000 50.2000 ;
	    RECT 76.4000 41.6000 77.2000 46.2000 ;
	    RECT 79.6000 41.6000 80.4000 49.8000 ;
	    RECT 82.8000 41.6000 83.6000 50.2000 ;
	    RECT 89.2000 41.6000 90.0000 49.0000 ;
	    RECT 92.4000 41.6000 93.2000 50.2000 ;
	    RECT 97.2000 41.6000 98.0000 50.2000 ;
	    RECT 0.4000 40.4000 102.0000 41.6000 ;
	    RECT 4.4000 31.8000 5.2000 40.4000 ;
	    RECT 6.0000 35.8000 6.8000 40.4000 ;
	    RECT 9.2000 32.2000 10.0000 40.4000 ;
	    RECT 15.6000 31.8000 16.4000 40.4000 ;
	    RECT 17.2000 35.8000 18.0000 40.4000 ;
	    RECT 20.4000 35.8000 21.2000 40.4000 ;
	    RECT 23.6000 35.8000 24.4000 40.4000 ;
	    RECT 26.8000 35.8000 27.6000 40.4000 ;
	    RECT 33.2000 35.8000 34.0000 40.4000 ;
	    RECT 36.4000 35.8000 37.2000 40.4000 ;
	    RECT 39.6000 35.8000 40.4000 40.4000 ;
	    RECT 41.2000 35.8000 42.0000 40.4000 ;
	    RECT 44.4000 35.8000 45.2000 40.4000 ;
	    RECT 47.6000 35.8000 48.4000 40.4000 ;
	    RECT 49.2000 35.8000 50.0000 40.4000 ;
	    RECT 52.4000 35.8000 53.2000 40.4000 ;
	    RECT 55.6000 32.2000 56.4000 40.4000 ;
	    RECT 58.8000 35.8000 59.6000 40.4000 ;
	    RECT 60.4000 35.8000 61.2000 40.4000 ;
	    RECT 63.6000 35.8000 64.4000 40.4000 ;
	    RECT 66.8000 35.8000 67.6000 40.4000 ;
	    RECT 68.4000 35.8000 69.2000 40.4000 ;
	    RECT 71.6000 35.8000 72.4000 40.4000 ;
	    RECT 78.0000 35.8000 78.8000 40.4000 ;
	    RECT 81.2000 35.8000 82.0000 40.4000 ;
	    RECT 84.4000 35.8000 85.2000 40.4000 ;
	    RECT 87.6000 35.8000 88.4000 40.4000 ;
	    RECT 92.4000 31.8000 93.2000 40.4000 ;
	    RECT 95.6000 32.2000 96.4000 40.4000 ;
	    RECT 98.8000 35.8000 99.6000 40.4000 ;
	    RECT 2.8000 1.6000 3.6000 9.0000 ;
	    RECT 6.0000 1.6000 6.8000 10.2000 ;
	    RECT 10.8000 1.6000 11.6000 10.2000 ;
	    RECT 15.6000 1.6000 16.4000 6.2000 ;
	    RECT 18.8000 1.6000 19.6000 9.8000 ;
	    RECT 23.6000 1.6000 24.4000 9.0000 ;
	    RECT 31.6000 1.6000 32.4000 10.2000 ;
	    RECT 38.0000 1.6000 38.8000 9.8000 ;
	    RECT 41.2000 1.6000 42.0000 6.2000 ;
	    RECT 46.0000 1.6000 46.8000 10.2000 ;
	    RECT 47.6000 1.6000 48.4000 10.2000 ;
	    RECT 55.6000 1.6000 56.4000 10.2000 ;
	    RECT 57.2000 1.6000 58.0000 6.2000 ;
	    RECT 60.4000 1.6000 61.2000 9.8000 ;
	    RECT 63.6000 1.6000 64.4000 6.2000 ;
	    RECT 66.8000 1.6000 67.6000 6.2000 ;
	    RECT 70.0000 1.6000 70.8000 9.0000 ;
	    RECT 79.6000 1.6000 80.4000 6.2000 ;
	    RECT 81.2000 1.6000 82.0000 10.2000 ;
	    RECT 86.0000 1.6000 86.8000 6.2000 ;
	    RECT 89.2000 1.6000 90.0000 9.8000 ;
	    RECT 95.6000 1.6000 96.4000 10.2000 ;
	    RECT 98.8000 1.6000 99.6000 9.0000 ;
	    RECT 0.4000 0.4000 102.0000 1.6000 ;
         LAYER metal2 ;
	    RECT 26.4000 80.6000 31.2000 81.4000 ;
	    RECT 26.4000 40.6000 31.2000 41.4000 ;
	    RECT 26.4000 0.6000 31.2000 1.4000 ;
         LAYER M3 ;
	    RECT 26.4000 80.4000 31.2000 81.6000 ;
	    RECT 26.4000 40.4000 31.2000 41.6000 ;
	    RECT 26.4000 0.4000 31.2000 1.6000 ;
         LAYER M4 ;
	    RECT 26.4000 -4.0000 31.2000 84.0000 ;
      END
   END vdd
   PIN gnd
      PORT
         LAYER M1 ;
	    RECT 1.2000 61.6000 2.0000 64.2000 ;
	    RECT 4.4000 61.6000 5.2000 64.2000 ;
	    RECT 8.6000 61.6000 9.4000 66.0000 ;
	    RECT 12.4000 61.6000 13.2000 64.2000 ;
	    RECT 15.6000 61.6000 16.4000 64.2000 ;
	    RECT 19.8000 61.6000 20.6000 66.0000 ;
	    RECT 23.6000 61.6000 24.4000 64.2000 ;
	    RECT 26.8000 61.6000 27.6000 64.2000 ;
	    RECT 33.2000 61.6000 34.0000 64.2000 ;
	    RECT 36.4000 61.6000 37.2000 64.2000 ;
	    RECT 39.6000 61.6000 40.4000 66.2000 ;
	    RECT 44.4000 61.6000 45.2000 66.2000 ;
	    RECT 47.6000 61.6000 48.4000 64.2000 ;
	    RECT 50.8000 61.6000 51.6000 64.2000 ;
	    RECT 54.6000 61.6000 55.4000 66.0000 ;
	    RECT 58.8000 61.6000 59.6000 64.2000 ;
	    RECT 62.0000 61.6000 62.8000 64.2000 ;
	    RECT 66.8000 61.6000 67.6000 66.2000 ;
	    RECT 70.0000 61.6000 70.8000 64.2000 ;
	    RECT 76.4000 61.6000 77.2000 64.2000 ;
	    RECT 79.6000 61.6000 80.4000 64.2000 ;
	    RECT 83.4000 61.6000 84.2000 66.0000 ;
	    RECT 87.6000 61.6000 88.4000 64.2000 ;
	    RECT 90.8000 61.6000 91.6000 64.2000 ;
	    RECT 94.6000 61.6000 95.4000 66.0000 ;
	    RECT 0.4000 60.4000 102.0000 61.6000 ;
	    RECT 1.2000 57.8000 2.0000 60.4000 ;
	    RECT 6.0000 57.8000 6.8000 60.4000 ;
	    RECT 7.6000 55.8000 8.4000 60.4000 ;
	    RECT 15.6000 55.8000 16.4000 60.4000 ;
	    RECT 17.2000 55.8000 18.0000 60.4000 ;
	    RECT 24.6000 56.0000 25.4000 60.4000 ;
	    RECT 36.4000 55.8000 37.2000 60.4000 ;
	    RECT 41.2000 55.8000 42.0000 60.4000 ;
	    RECT 44.4000 57.8000 45.2000 60.4000 ;
	    RECT 49.2000 55.8000 50.0000 60.4000 ;
	    RECT 52.4000 57.8000 53.2000 60.4000 ;
	    RECT 57.2000 55.8000 58.0000 60.4000 ;
	    RECT 60.4000 57.8000 61.2000 60.4000 ;
	    RECT 62.0000 57.8000 62.8000 60.4000 ;
	    RECT 65.2000 57.8000 66.0000 60.4000 ;
	    RECT 66.8000 57.8000 67.6000 60.4000 ;
	    RECT 70.0000 57.8000 70.8000 60.4000 ;
	    RECT 79.0000 56.0000 79.8000 60.4000 ;
	    RECT 82.8000 57.8000 83.6000 60.4000 ;
	    RECT 86.0000 57.8000 86.8000 60.4000 ;
	    RECT 89.2000 55.8000 90.0000 60.4000 ;
	    RECT 92.4000 57.8000 93.2000 60.4000 ;
	    RECT 95.6000 57.8000 96.4000 60.4000 ;
	    RECT 97.2000 57.8000 98.0000 60.4000 ;
	    RECT 100.4000 57.8000 101.2000 60.4000 ;
	    RECT 1.2000 21.6000 2.0000 24.2000 ;
	    RECT 4.4000 21.6000 5.2000 24.2000 ;
	    RECT 8.6000 21.6000 9.4000 26.0000 ;
	    RECT 12.4000 21.6000 13.2000 24.2000 ;
	    RECT 15.6000 21.6000 16.4000 24.2000 ;
	    RECT 17.2000 21.6000 18.0000 24.2000 ;
	    RECT 20.4000 21.6000 21.2000 24.2000 ;
	    RECT 23.6000 21.6000 24.4000 26.2000 ;
	    RECT 33.2000 21.6000 34.0000 24.2000 ;
	    RECT 36.4000 21.6000 37.2000 26.2000 ;
	    RECT 41.2000 21.6000 42.0000 26.2000 ;
	    RECT 47.6000 21.6000 48.4000 24.2000 ;
	    RECT 49.2000 21.6000 50.0000 26.2000 ;
	    RECT 56.2000 21.6000 57.0000 26.0000 ;
	    RECT 63.6000 21.6000 64.4000 26.2000 ;
	    RECT 66.8000 21.6000 67.6000 24.2000 ;
	    RECT 68.4000 21.6000 69.2000 26.2000 ;
	    RECT 81.2000 21.6000 82.0000 26.2000 ;
	    RECT 84.4000 21.6000 85.2000 24.2000 ;
	    RECT 87.6000 21.6000 88.4000 24.2000 ;
	    RECT 89.2000 21.6000 90.0000 24.2000 ;
	    RECT 92.4000 21.6000 93.2000 24.2000 ;
	    RECT 96.2000 21.6000 97.0000 26.0000 ;
	    RECT 0.4000 20.4000 102.0000 21.6000 ;
	    RECT 2.8000 15.8000 3.6000 20.4000 ;
	    RECT 6.0000 17.8000 6.8000 20.4000 ;
	    RECT 9.2000 17.8000 10.0000 20.4000 ;
	    RECT 10.8000 17.8000 11.6000 20.4000 ;
	    RECT 14.0000 17.8000 14.8000 20.4000 ;
	    RECT 18.2000 16.0000 19.0000 20.4000 ;
	    RECT 23.6000 15.8000 24.4000 20.4000 ;
	    RECT 31.6000 17.8000 32.4000 20.4000 ;
	    RECT 34.8000 17.8000 35.6000 20.4000 ;
	    RECT 38.6000 16.0000 39.4000 20.4000 ;
	    RECT 42.8000 17.8000 43.6000 20.4000 ;
	    RECT 46.0000 17.8000 46.8000 20.4000 ;
	    RECT 47.6000 17.8000 48.4000 20.4000 ;
	    RECT 50.8000 17.8000 51.6000 20.4000 ;
	    RECT 52.4000 17.8000 53.2000 20.4000 ;
	    RECT 55.6000 17.8000 56.4000 20.4000 ;
	    RECT 59.8000 16.0000 60.6000 20.4000 ;
	    RECT 66.8000 15.8000 67.6000 20.4000 ;
	    RECT 70.0000 15.8000 70.8000 20.4000 ;
	    RECT 79.6000 17.8000 80.4000 20.4000 ;
	    RECT 81.2000 17.8000 82.0000 20.4000 ;
	    RECT 84.4000 17.8000 85.2000 20.4000 ;
	    RECT 88.6000 16.0000 89.4000 20.4000 ;
	    RECT 92.4000 17.8000 93.2000 20.4000 ;
	    RECT 95.6000 17.8000 96.4000 20.4000 ;
	    RECT 98.8000 15.8000 99.6000 20.4000 ;
         LAYER metal2 ;
	    RECT 71.2000 60.6000 76.0000 61.4000 ;
	    RECT 71.2000 20.6000 76.0000 21.4000 ;
         LAYER M3 ;
	    RECT 71.2000 60.4000 76.0000 61.6000 ;
	    RECT 71.2000 20.4000 76.0000 21.6000 ;
         LAYER M4 ;
	    RECT 71.2000 -4.0000 76.0000 84.0000 ;
      END
   END gnd
   PIN sum_comp_1[0]
      PORT
         LAYER M1 ;
	    RECT 84.4000 69.6000 85.2000 70.4000 ;
	    RECT 90.8000 69.6000 91.6000 71.2000 ;
	    RECT 84.4000 68.8000 85.0000 69.6000 ;
	    RECT 84.0000 68.2000 85.0000 68.8000 ;
	    RECT 84.0000 68.0000 84.8000 68.2000 ;
         LAYER metal2 ;
	    RECT 89.3000 70.4000 89.9000 84.3000 ;
	    RECT 84.4000 69.6000 85.2000 70.4000 ;
	    RECT 89.2000 69.6000 90.0000 70.4000 ;
	    RECT 90.8000 69.6000 91.6000 70.4000 ;
         LAYER M3 ;
	    RECT 84.4000 70.3000 85.2000 70.4000 ;
	    RECT 89.2000 70.3000 90.0000 70.4000 ;
	    RECT 90.8000 70.3000 91.6000 70.4000 ;
	    RECT 84.4000 69.7000 91.6000 70.3000 ;
	    RECT 84.4000 69.6000 85.2000 69.7000 ;
	    RECT 89.2000 69.6000 90.0000 69.7000 ;
	    RECT 90.8000 69.6000 91.6000 69.7000 ;
      END
   END sum_comp_1[0]
   PIN sum_comp_1[1]
      PORT
         LAYER M1 ;
	    RECT 95.6000 69.6000 96.4000 70.4000 ;
	    RECT 95.6000 68.8000 96.2000 69.6000 ;
	    RECT 95.2000 68.2000 96.2000 68.8000 ;
	    RECT 95.2000 68.0000 96.0000 68.2000 ;
	    RECT 95.6000 50.8000 96.4000 52.4000 ;
         LAYER metal2 ;
	    RECT 95.6000 69.6000 96.4000 70.4000 ;
	    RECT 95.7000 52.4000 96.3000 69.6000 ;
	    RECT 95.6000 51.6000 96.4000 52.4000 ;
         LAYER M3 ;
	    RECT 95.6000 52.3000 96.4000 52.4000 ;
	    RECT 95.6000 51.7000 104.3000 52.3000 ;
	    RECT 95.6000 51.6000 96.4000 51.7000 ;
      END
   END sum_comp_1[1]
   PIN sum_comp_1[2]
      PORT
         LAYER M1 ;
	    RECT 1.2000 69.6000 2.0000 71.2000 ;
	    RECT 7.6000 69.6000 8.4000 70.4000 ;
	    RECT 7.8000 68.8000 8.4000 69.6000 ;
	    RECT 7.8000 68.2000 8.8000 68.8000 ;
	    RECT 8.0000 68.0000 8.8000 68.2000 ;
         LAYER metal2 ;
	    RECT 1.2000 69.6000 2.0000 70.4000 ;
	    RECT 7.6000 69.6000 8.4000 70.4000 ;
         LAYER M3 ;
	    RECT 1.2000 70.3000 2.0000 70.4000 ;
	    RECT 7.6000 70.3000 8.4000 70.4000 ;
	    RECT -1.9000 69.7000 8.4000 70.3000 ;
	    RECT 1.2000 69.6000 2.0000 69.7000 ;
	    RECT 7.6000 69.6000 8.4000 69.7000 ;
      END
   END sum_comp_1[2]
   PIN sum_comp_1[3]
      PORT
         LAYER M1 ;
	    RECT 1.2000 29.6000 2.0000 31.2000 ;
	    RECT 7.6000 29.6000 8.4000 30.4000 ;
	    RECT 7.8000 28.8000 8.4000 29.6000 ;
	    RECT 7.8000 28.2000 8.8000 28.8000 ;
	    RECT 8.0000 28.0000 8.8000 28.2000 ;
         LAYER metal2 ;
	    RECT 1.2000 31.6000 2.0000 32.4000 ;
	    RECT 7.6000 31.6000 8.4000 32.4000 ;
	    RECT 1.3000 30.4000 1.9000 31.6000 ;
	    RECT 7.7000 30.4000 8.3000 31.6000 ;
	    RECT 1.2000 29.6000 2.0000 30.4000 ;
	    RECT 7.6000 29.6000 8.4000 30.4000 ;
         LAYER M3 ;
	    RECT 1.2000 32.3000 2.0000 32.4000 ;
	    RECT 7.6000 32.3000 8.4000 32.4000 ;
	    RECT -1.9000 31.7000 8.4000 32.3000 ;
	    RECT 1.2000 31.6000 2.0000 31.7000 ;
	    RECT 7.6000 31.6000 8.4000 31.7000 ;
      END
   END sum_comp_1[3]
   PIN sum_comp_1[4]
      PORT
         LAYER M1 ;
	    RECT 59.2000 13.8000 60.0000 14.0000 ;
	    RECT 59.0000 13.2000 60.0000 13.8000 ;
	    RECT 59.0000 12.4000 59.6000 13.2000 ;
	    RECT 52.4000 10.8000 53.2000 12.4000 ;
	    RECT 58.8000 11.6000 59.6000 12.4000 ;
         LAYER metal2 ;
	    RECT 52.4000 11.6000 53.2000 12.4000 ;
	    RECT 54.0000 11.6000 54.8000 12.4000 ;
	    RECT 58.8000 11.6000 59.6000 12.4000 ;
	    RECT 54.1000 -2.3000 54.7000 11.6000 ;
         LAYER M3 ;
	    RECT 52.4000 12.3000 53.2000 12.4000 ;
	    RECT 54.0000 12.3000 54.8000 12.4000 ;
	    RECT 58.8000 12.3000 59.6000 12.4000 ;
	    RECT 52.4000 11.7000 59.6000 12.3000 ;
	    RECT 52.4000 11.6000 53.2000 11.7000 ;
	    RECT 54.0000 11.6000 54.8000 11.7000 ;
	    RECT 58.8000 11.6000 59.6000 11.7000 ;
      END
   END sum_comp_1[4]
   PIN sum_comp_1[5]
      PORT
         LAYER M1 ;
	    RECT 100.4000 50.8000 101.2000 52.4000 ;
	    RECT 97.2000 29.6000 98.0000 30.4000 ;
	    RECT 97.2000 28.8000 97.8000 29.6000 ;
	    RECT 96.8000 28.2000 97.8000 28.8000 ;
	    RECT 96.8000 28.0000 97.6000 28.2000 ;
         LAYER metal2 ;
	    RECT 100.4000 51.6000 101.2000 52.4000 ;
	    RECT 100.5000 50.4000 101.1000 51.6000 ;
	    RECT 100.4000 49.6000 101.2000 50.4000 ;
	    RECT 97.2000 29.6000 98.0000 30.4000 ;
         LAYER M3 ;
	    RECT 100.4000 64.3000 101.2000 64.4000 ;
	    RECT 100.4000 63.7000 104.3000 64.3000 ;
	    RECT 100.4000 63.6000 101.2000 63.7000 ;
	    RECT 100.4000 49.6000 101.2000 50.4000 ;
	    RECT 97.2000 30.3000 98.0000 30.4000 ;
	    RECT 100.4000 30.3000 101.2000 30.4000 ;
	    RECT 97.2000 29.7000 101.2000 30.3000 ;
	    RECT 97.2000 29.6000 98.0000 29.7000 ;
	    RECT 100.4000 29.6000 101.2000 29.7000 ;
         LAYER M4 ;
	    RECT 100.2000 29.4000 101.4000 64.6000 ;
      END
   END sum_comp_1[5]
   PIN sum_comp_2[0]
      PORT
         LAYER M1 ;
	    RECT 86.0000 68.3000 86.8000 70.4000 ;
	    RECT 86.0000 67.7000 88.3000 68.3000 ;
	    RECT 86.0000 67.6000 86.8000 67.7000 ;
	    RECT 87.7000 66.4000 88.3000 67.7000 ;
	    RECT 87.6000 64.8000 88.4000 66.4000 ;
         LAYER metal2 ;
	    RECT 82.9000 80.4000 83.5000 84.3000 ;
	    RECT 82.8000 79.6000 83.6000 80.4000 ;
	    RECT 86.0000 79.6000 86.8000 80.4000 ;
	    RECT 86.1000 70.4000 86.7000 79.6000 ;
	    RECT 86.0000 69.6000 86.8000 70.4000 ;
         LAYER M3 ;
	    RECT 82.8000 80.3000 83.6000 80.4000 ;
	    RECT 86.0000 80.3000 86.8000 80.4000 ;
	    RECT 82.8000 79.7000 86.8000 80.3000 ;
	    RECT 82.8000 79.6000 83.6000 79.7000 ;
	    RECT 86.0000 79.6000 86.8000 79.7000 ;
      END
   END sum_comp_2[0]
   PIN sum_comp_2[1]
      PORT
         LAYER M1 ;
	    RECT 97.2000 68.3000 98.0000 69.2000 ;
	    RECT 100.4000 68.3000 101.2000 68.4000 ;
	    RECT 97.2000 67.7000 101.2000 68.3000 ;
	    RECT 97.2000 67.6000 98.0000 67.7000 ;
	    RECT 100.4000 67.6000 101.2000 67.7000 ;
	    RECT 92.4000 55.6000 93.2000 57.2000 ;
         LAYER metal2 ;
	    RECT 100.4000 67.6000 101.2000 68.4000 ;
	    RECT 100.5000 60.4000 101.1000 67.6000 ;
	    RECT 92.4000 59.6000 93.2000 60.4000 ;
	    RECT 100.4000 59.6000 101.2000 60.4000 ;
	    RECT 92.5000 56.4000 93.1000 59.6000 ;
	    RECT 92.4000 55.6000 93.2000 56.4000 ;
         LAYER M3 ;
	    RECT 92.4000 60.3000 93.2000 60.4000 ;
	    RECT 100.4000 60.3000 101.2000 60.4000 ;
	    RECT 92.4000 59.7000 104.3000 60.3000 ;
	    RECT 92.4000 59.6000 93.2000 59.7000 ;
	    RECT 100.4000 59.6000 101.2000 59.7000 ;
      END
   END sum_comp_2[1]
   PIN sum_comp_2[2]
      PORT
         LAYER M1 ;
	    RECT 6.0000 68.3000 6.8000 69.2000 ;
	    RECT 4.5000 67.7000 6.8000 68.3000 ;
	    RECT 4.5000 66.4000 5.1000 67.7000 ;
	    RECT 6.0000 67.6000 6.8000 67.7000 ;
	    RECT 4.4000 64.8000 5.2000 66.4000 ;
         LAYER metal2 ;
	    RECT 4.4000 65.6000 5.2000 66.4000 ;
         LAYER M3 ;
	    RECT 4.4000 66.3000 5.2000 66.4000 ;
	    RECT -1.9000 65.7000 5.2000 66.3000 ;
	    RECT 4.4000 65.6000 5.2000 65.7000 ;
      END
   END sum_comp_2[2]
   PIN sum_comp_2[3]
      PORT
         LAYER M1 ;
	    RECT 4.4000 28.3000 5.2000 28.4000 ;
	    RECT 6.0000 28.3000 6.8000 29.2000 ;
	    RECT 4.4000 27.7000 6.8000 28.3000 ;
	    RECT 4.4000 27.6000 5.2000 27.7000 ;
	    RECT 6.0000 27.6000 6.8000 27.7000 ;
	    RECT 4.5000 26.4000 5.1000 27.6000 ;
	    RECT 4.4000 24.8000 5.2000 26.4000 ;
         LAYER metal2 ;
	    RECT 4.4000 27.6000 5.2000 28.4000 ;
         LAYER M3 ;
	    RECT 4.4000 28.3000 5.2000 28.4000 ;
	    RECT -1.9000 27.7000 5.2000 28.3000 ;
	    RECT 4.4000 27.6000 5.2000 27.7000 ;
      END
   END sum_comp_2[3]
   PIN sum_comp_2[4]
      PORT
         LAYER M1 ;
	    RECT 55.6000 15.6000 56.4000 17.2000 ;
	    RECT 55.7000 14.3000 56.3000 15.6000 ;
	    RECT 57.2000 14.3000 58.0000 14.4000 ;
	    RECT 55.7000 13.7000 58.0000 14.3000 ;
	    RECT 57.2000 11.6000 58.0000 13.7000 ;
         LAYER metal2 ;
	    RECT 57.2000 11.6000 58.0000 12.4000 ;
	    RECT 57.3000 -2.3000 57.9000 11.6000 ;
      END
   END sum_comp_2[4]
   PIN sum_comp_2[5]
      PORT
         LAYER M1 ;
	    RECT 97.2000 55.6000 98.0000 57.2000 ;
	    RECT 100.4000 30.3000 101.2000 30.4000 ;
	    RECT 98.8000 29.7000 101.2000 30.3000 ;
	    RECT 98.8000 27.6000 99.6000 29.7000 ;
	    RECT 100.4000 29.6000 101.2000 29.7000 ;
         LAYER metal2 ;
	    RECT 97.2000 55.6000 98.0000 56.4000 ;
	    RECT 97.3000 32.4000 97.9000 55.6000 ;
	    RECT 97.2000 31.6000 98.0000 32.4000 ;
	    RECT 100.4000 31.6000 101.2000 32.4000 ;
	    RECT 100.5000 30.4000 101.1000 31.6000 ;
	    RECT 100.4000 29.6000 101.2000 30.4000 ;
         LAYER M3 ;
	    RECT 97.2000 32.3000 98.0000 32.4000 ;
	    RECT 100.4000 32.3000 101.2000 32.4000 ;
	    RECT 97.2000 31.7000 104.3000 32.3000 ;
	    RECT 97.2000 31.6000 98.0000 31.7000 ;
	    RECT 100.4000 31.6000 101.2000 31.7000 ;
      END
   END sum_comp_2[5]
   PIN c_in
      PORT
         LAYER M1 ;
	    RECT 63.6000 71.6000 64.4000 74.4000 ;
	    RECT 57.2000 68.3000 58.0000 69.2000 ;
	    RECT 58.8000 68.3000 59.6000 68.4000 ;
	    RECT 57.2000 67.7000 59.6000 68.3000 ;
	    RECT 57.2000 67.6000 58.0000 67.7000 ;
	    RECT 58.8000 67.6000 59.6000 67.7000 ;
	    RECT 58.8000 64.8000 59.6000 66.4000 ;
         LAYER metal2 ;
	    RECT 63.7000 74.4000 64.3000 84.3000 ;
	    RECT 63.6000 73.6000 64.4000 74.4000 ;
	    RECT 63.7000 70.4000 64.3000 73.6000 ;
	    RECT 58.8000 69.6000 59.6000 70.4000 ;
	    RECT 63.6000 69.6000 64.4000 70.4000 ;
	    RECT 58.9000 68.4000 59.5000 69.6000 ;
	    RECT 58.8000 67.6000 59.6000 68.4000 ;
	    RECT 58.9000 66.4000 59.5000 67.6000 ;
	    RECT 58.8000 65.6000 59.6000 66.4000 ;
         LAYER M3 ;
	    RECT 58.8000 70.3000 59.6000 70.4000 ;
	    RECT 63.6000 70.3000 64.4000 70.4000 ;
	    RECT 58.8000 69.7000 64.4000 70.3000 ;
	    RECT 58.8000 69.6000 59.6000 69.7000 ;
	    RECT 63.6000 69.6000 64.4000 69.7000 ;
      END
   END c_in
   PIN result[0]
      PORT
         LAYER M1 ;
	    RECT 42.8000 71.8000 43.6000 79.8000 ;
	    RECT 42.8000 69.6000 43.4000 71.8000 ;
	    RECT 42.8000 62.2000 43.6000 69.6000 ;
         LAYER metal2 ;
	    RECT 42.9000 83.7000 45.1000 84.3000 ;
	    RECT 42.9000 78.4000 43.5000 83.7000 ;
	    RECT 42.8000 77.6000 43.6000 78.4000 ;
      END
   END result[0]
   PIN result[1]
      PORT
         LAYER M1 ;
	    RECT 90.8000 52.4000 91.6000 59.8000 ;
	    RECT 91.0000 50.2000 91.6000 52.4000 ;
	    RECT 90.8000 42.2000 91.6000 50.2000 ;
         LAYER metal2 ;
	    RECT 90.8000 57.6000 91.6000 58.4000 ;
         LAYER M3 ;
	    RECT 90.8000 58.3000 91.6000 58.4000 ;
	    RECT 90.8000 57.7000 102.7000 58.3000 ;
	    RECT 90.8000 57.6000 91.6000 57.7000 ;
	    RECT 102.1000 56.3000 102.7000 57.7000 ;
	    RECT 102.1000 55.7000 104.3000 56.3000 ;
      END
   END result[1]
   PIN result[2]
      PORT
         LAYER M1 ;
	    RECT 41.2000 71.8000 42.0000 79.8000 ;
	    RECT 41.4000 69.6000 42.0000 71.8000 ;
	    RECT 41.2000 62.2000 42.0000 69.6000 ;
         LAYER metal2 ;
	    RECT 39.7000 83.7000 41.9000 84.3000 ;
	    RECT 41.3000 78.4000 41.9000 83.7000 ;
	    RECT 41.2000 77.6000 42.0000 78.4000 ;
      END
   END result[2]
   PIN result[3]
      PORT
         LAYER M1 ;
	    RECT 1.2000 12.4000 2.0000 19.8000 ;
	    RECT 1.2000 10.2000 1.8000 12.4000 ;
	    RECT 1.2000 2.2000 2.0000 10.2000 ;
         LAYER metal2 ;
	    RECT 1.2000 9.6000 2.0000 10.4000 ;
	    RECT 1.3000 8.4000 1.9000 9.6000 ;
	    RECT 1.2000 7.6000 2.0000 8.4000 ;
         LAYER M3 ;
	    RECT 1.2000 10.3000 2.0000 10.4000 ;
	    RECT -1.9000 9.7000 2.0000 10.3000 ;
	    RECT 1.2000 9.6000 2.0000 9.7000 ;
      END
   END result[3]
   PIN result[4]
      PORT
         LAYER M1 ;
	    RECT 22.0000 12.4000 22.8000 19.8000 ;
	    RECT 22.0000 10.2000 22.6000 12.4000 ;
	    RECT 22.0000 2.2000 22.8000 10.2000 ;
         LAYER metal2 ;
	    RECT 22.0000 3.6000 22.8000 4.4000 ;
	    RECT 22.1000 -1.7000 22.7000 3.6000 ;
	    RECT 22.1000 -2.3000 24.3000 -1.7000 ;
      END
   END result[4]
   PIN result[5]
      PORT
         LAYER M1 ;
	    RECT 100.4000 12.4000 101.2000 19.8000 ;
	    RECT 100.6000 10.2000 101.2000 12.4000 ;
	    RECT 100.4000 2.2000 101.2000 10.2000 ;
         LAYER metal2 ;
	    RECT 100.4000 9.6000 101.2000 10.4000 ;
	    RECT 100.5000 8.4000 101.1000 9.6000 ;
	    RECT 100.4000 7.6000 101.2000 8.4000 ;
         LAYER M3 ;
	    RECT 100.4000 10.3000 101.2000 10.4000 ;
	    RECT 100.4000 9.7000 104.3000 10.3000 ;
	    RECT 100.4000 9.6000 101.2000 9.7000 ;
      END
   END result[5]
   PIN c_out
      PORT
         LAYER M1 ;
	    RECT 71.6000 12.4000 72.4000 19.8000 ;
	    RECT 71.8000 10.2000 72.4000 12.4000 ;
	    RECT 71.6000 4.3000 72.4000 10.2000 ;
	    RECT 76.4000 4.3000 77.2000 4.4000 ;
	    RECT 71.6000 3.7000 77.2000 4.3000 ;
	    RECT 71.6000 2.2000 72.4000 3.7000 ;
	    RECT 76.4000 3.6000 77.2000 3.7000 ;
         LAYER metal2 ;
	    RECT 76.4000 3.6000 77.2000 4.4000 ;
	    RECT 76.5000 -2.3000 77.1000 3.6000 ;
      END
   END c_out
   OBS
         LAYER M1 ;
	    RECT 1.8000 72.6000 2.6000 79.8000 ;
	    RECT 7.6000 75.8000 8.4000 79.8000 ;
	    RECT 1.8000 71.8000 3.6000 72.6000 ;
	    RECT 2.8000 68.4000 3.4000 71.8000 ;
	    RECT 7.8000 71.6000 8.4000 75.8000 ;
	    RECT 10.8000 71.8000 11.6000 79.8000 ;
	    RECT 15.0000 74.3000 15.8000 79.8000 ;
	    RECT 18.8000 75.8000 19.6000 79.8000 ;
	    RECT 17.2000 74.3000 18.0000 74.4000 ;
	    RECT 15.0000 73.7000 18.0000 74.3000 ;
	    RECT 15.0000 72.6000 15.8000 73.7000 ;
	    RECT 17.2000 73.6000 18.0000 73.7000 ;
	    RECT 14.0000 71.8000 15.8000 72.6000 ;
	    RECT 7.8000 71.0000 10.2000 71.6000 ;
	    RECT 2.8000 67.6000 3.6000 68.4000 ;
	    RECT 9.6000 67.6000 10.2000 71.0000 ;
	    RECT 11.0000 70.4000 11.6000 71.8000 ;
	    RECT 10.8000 70.3000 11.6000 70.4000 ;
	    RECT 12.4000 70.3000 13.2000 70.4000 ;
	    RECT 10.8000 69.7000 13.2000 70.3000 ;
	    RECT 10.8000 69.6000 11.6000 69.7000 ;
	    RECT 12.4000 69.6000 13.2000 69.7000 ;
	    RECT 1.2000 66.3000 2.0000 66.4000 ;
	    RECT 2.8000 66.3000 3.4000 67.6000 ;
	    RECT 9.6000 67.4000 10.4000 67.6000 ;
	    RECT 7.4000 67.0000 10.4000 67.4000 ;
	    RECT 6.2000 66.8000 10.4000 67.0000 ;
	    RECT 6.2000 66.4000 8.0000 66.8000 ;
	    RECT 1.2000 65.7000 3.5000 66.3000 ;
	    RECT 6.2000 66.2000 6.8000 66.4000 ;
	    RECT 11.0000 66.2000 11.6000 69.6000 ;
	    RECT 14.2000 68.4000 14.8000 71.8000 ;
	    RECT 19.0000 71.6000 19.6000 75.8000 ;
	    RECT 22.0000 71.6000 22.8000 79.8000 ;
	    RECT 24.2000 72.6000 25.0000 79.8000 ;
	    RECT 33.8000 72.6000 34.6000 79.8000 ;
	    RECT 24.2000 71.8000 26.0000 72.6000 ;
	    RECT 33.8000 71.8000 35.6000 72.6000 ;
	    RECT 38.0000 72.4000 38.8000 79.8000 ;
	    RECT 46.0000 72.4000 46.8000 79.8000 ;
	    RECT 48.2000 74.4000 49.0000 79.8000 ;
	    RECT 47.6000 73.6000 49.0000 74.4000 ;
	    RECT 38.0000 71.8000 40.2000 72.4000 ;
	    RECT 15.6000 69.6000 16.4000 71.2000 ;
	    RECT 19.0000 71.0000 21.4000 71.6000 ;
	    RECT 18.8000 69.6000 19.6000 70.4000 ;
	    RECT 14.0000 67.6000 14.8000 68.4000 ;
	    RECT 17.2000 67.6000 18.0000 69.2000 ;
	    RECT 19.0000 68.8000 19.6000 69.6000 ;
	    RECT 19.0000 68.2000 20.0000 68.8000 ;
	    RECT 19.2000 68.0000 20.0000 68.2000 ;
	    RECT 20.8000 67.6000 21.4000 71.0000 ;
	    RECT 22.2000 70.4000 22.8000 71.6000 ;
	    RECT 22.0000 69.6000 22.8000 70.4000 ;
	    RECT 23.6000 69.6000 24.4000 71.2000 ;
	    RECT 1.2000 65.6000 2.0000 65.7000 ;
	    RECT 2.8000 64.2000 3.4000 65.7000 ;
	    RECT 2.8000 62.2000 3.6000 64.2000 ;
	    RECT 6.0000 62.2000 6.8000 66.2000 ;
	    RECT 10.2000 65.2000 11.6000 66.2000 ;
	    RECT 10.2000 62.2000 11.0000 65.2000 ;
	    RECT 12.4000 64.8000 13.2000 66.4000 ;
	    RECT 14.2000 64.2000 14.8000 67.6000 ;
	    RECT 20.8000 67.4000 21.6000 67.6000 ;
	    RECT 18.6000 67.0000 21.6000 67.4000 ;
	    RECT 17.4000 66.8000 21.6000 67.0000 ;
	    RECT 17.4000 66.4000 19.2000 66.8000 ;
	    RECT 17.4000 66.2000 18.0000 66.4000 ;
	    RECT 22.2000 66.2000 22.8000 69.6000 ;
	    RECT 14.0000 62.2000 14.8000 64.2000 ;
	    RECT 17.2000 62.2000 18.0000 66.2000 ;
	    RECT 21.4000 65.2000 22.8000 66.2000 ;
	    RECT 25.2000 68.4000 25.8000 71.8000 ;
	    RECT 33.2000 69.6000 34.0000 71.2000 ;
	    RECT 34.8000 70.3000 35.4000 71.8000 ;
	    RECT 39.6000 71.2000 40.2000 71.8000 ;
	    RECT 44.6000 71.8000 46.8000 72.4000 ;
	    RECT 48.2000 72.6000 49.0000 73.6000 ;
	    RECT 48.2000 71.8000 50.0000 72.6000 ;
	    RECT 52.4000 71.8000 53.2000 79.8000 ;
	    RECT 55.6000 75.8000 56.4000 79.8000 ;
	    RECT 44.6000 71.2000 45.2000 71.8000 ;
	    RECT 39.6000 70.4000 40.8000 71.2000 ;
	    RECT 44.0000 70.4000 45.2000 71.2000 ;
	    RECT 38.0000 70.3000 38.8000 70.4000 ;
	    RECT 34.8000 69.7000 38.8000 70.3000 ;
	    RECT 34.8000 68.4000 35.4000 69.7000 ;
	    RECT 38.0000 68.8000 38.8000 69.7000 ;
	    RECT 25.2000 67.6000 26.0000 68.4000 ;
	    RECT 34.8000 67.6000 35.6000 68.4000 ;
	    RECT 25.2000 66.4000 25.8000 67.6000 ;
	    RECT 25.2000 65.6000 26.0000 66.4000 ;
	    RECT 21.4000 62.2000 22.2000 65.2000 ;
	    RECT 25.2000 64.2000 25.8000 65.6000 ;
	    RECT 26.8000 64.8000 27.6000 66.4000 ;
	    RECT 34.8000 64.2000 35.4000 67.6000 ;
	    RECT 39.6000 67.4000 40.2000 70.4000 ;
	    RECT 38.0000 66.8000 40.2000 67.4000 ;
	    RECT 44.6000 67.4000 45.2000 70.4000 ;
	    RECT 46.0000 68.8000 46.8000 70.4000 ;
	    RECT 47.6000 69.6000 48.4000 71.2000 ;
	    RECT 49.2000 68.4000 49.8000 71.8000 ;
	    RECT 52.4000 70.4000 53.0000 71.8000 ;
	    RECT 55.6000 71.6000 56.2000 75.8000 ;
	    RECT 61.4000 72.6000 62.2000 79.8000 ;
	    RECT 60.4000 71.8000 62.2000 72.6000 ;
	    RECT 53.8000 71.0000 56.2000 71.6000 ;
	    RECT 50.8000 70.3000 51.6000 70.4000 ;
	    RECT 52.4000 70.3000 53.2000 70.4000 ;
	    RECT 50.8000 69.7000 53.2000 70.3000 ;
	    RECT 50.8000 69.6000 51.6000 69.7000 ;
	    RECT 52.4000 69.6000 53.2000 69.7000 ;
	    RECT 49.2000 67.6000 50.0000 68.4000 ;
	    RECT 44.6000 66.8000 46.8000 67.4000 ;
	    RECT 36.4000 64.8000 37.2000 66.4000 ;
	    RECT 25.2000 62.2000 26.0000 64.2000 ;
	    RECT 34.8000 62.2000 35.6000 64.2000 ;
	    RECT 38.0000 62.2000 38.8000 66.8000 ;
	    RECT 46.0000 62.2000 46.8000 66.8000 ;
	    RECT 49.2000 64.2000 49.8000 67.6000 ;
	    RECT 50.8000 64.8000 51.6000 66.4000 ;
	    RECT 52.4000 66.2000 53.0000 69.6000 ;
	    RECT 53.8000 67.6000 54.4000 71.0000 ;
	    RECT 55.6000 69.6000 56.4000 70.4000 ;
	    RECT 55.6000 68.8000 56.2000 69.6000 ;
	    RECT 55.2000 68.2000 56.2000 68.8000 ;
	    RECT 60.6000 68.4000 61.2000 71.8000 ;
	    RECT 62.0000 69.6000 62.8000 71.2000 ;
	    RECT 55.2000 68.0000 56.0000 68.2000 ;
	    RECT 60.4000 67.6000 61.2000 68.4000 ;
	    RECT 53.6000 67.4000 54.4000 67.6000 ;
	    RECT 53.6000 67.0000 56.6000 67.4000 ;
	    RECT 53.6000 66.8000 57.8000 67.0000 ;
	    RECT 56.0000 66.4000 57.8000 66.8000 ;
	    RECT 60.6000 66.4000 61.2000 67.6000 ;
	    RECT 57.2000 66.2000 57.8000 66.4000 ;
	    RECT 52.4000 65.2000 53.8000 66.2000 ;
	    RECT 49.2000 62.2000 50.0000 64.2000 ;
	    RECT 53.0000 62.2000 53.8000 65.2000 ;
	    RECT 57.2000 62.2000 58.0000 66.2000 ;
	    RECT 60.4000 65.6000 61.2000 66.4000 ;
	    RECT 65.2000 66.2000 66.0000 79.8000 ;
	    RECT 66.8000 68.3000 67.6000 68.4000 ;
	    RECT 68.4000 68.3000 69.2000 79.8000 ;
	    RECT 77.0000 72.6000 77.8000 79.8000 ;
	    RECT 77.0000 71.8000 78.8000 72.6000 ;
	    RECT 78.0000 71.6000 78.8000 71.8000 ;
	    RECT 81.2000 71.8000 82.0000 79.8000 ;
	    RECT 84.4000 75.8000 85.2000 79.8000 ;
	    RECT 76.4000 69.6000 77.2000 71.2000 ;
	    RECT 66.8000 67.7000 69.2000 68.3000 ;
	    RECT 66.8000 66.8000 67.6000 67.7000 ;
	    RECT 60.6000 64.2000 61.2000 65.6000 ;
	    RECT 64.2000 65.6000 66.0000 66.2000 ;
	    RECT 64.2000 64.4000 65.0000 65.6000 ;
	    RECT 60.4000 62.2000 61.2000 64.2000 ;
	    RECT 63.6000 63.6000 65.0000 64.4000 ;
	    RECT 64.2000 62.2000 65.0000 63.6000 ;
	    RECT 68.4000 62.2000 69.2000 67.7000 ;
	    RECT 78.0000 68.4000 78.6000 71.6000 ;
	    RECT 81.2000 70.4000 81.8000 71.8000 ;
	    RECT 84.4000 71.6000 85.0000 75.8000 ;
	    RECT 90.2000 72.6000 91.0000 79.8000 ;
	    RECT 89.2000 71.8000 91.0000 72.6000 ;
	    RECT 92.4000 71.8000 93.2000 79.8000 ;
	    RECT 95.6000 75.8000 96.4000 79.8000 ;
	    RECT 82.6000 71.0000 85.0000 71.6000 ;
	    RECT 81.2000 69.6000 82.0000 70.4000 ;
	    RECT 78.0000 67.6000 78.8000 68.4000 ;
	    RECT 70.0000 64.8000 70.8000 66.4000 ;
	    RECT 78.0000 64.2000 78.6000 67.6000 ;
	    RECT 79.6000 64.8000 80.4000 66.4000 ;
	    RECT 81.2000 66.2000 81.8000 69.6000 ;
	    RECT 82.6000 67.6000 83.2000 71.0000 ;
	    RECT 89.4000 68.4000 90.0000 71.8000 ;
	    RECT 89.2000 67.6000 90.0000 68.4000 ;
	    RECT 82.4000 67.4000 83.2000 67.6000 ;
	    RECT 82.4000 67.0000 85.4000 67.4000 ;
	    RECT 82.4000 66.8000 86.6000 67.0000 ;
	    RECT 84.8000 66.4000 86.6000 66.8000 ;
	    RECT 89.4000 66.4000 90.0000 67.6000 ;
	    RECT 86.0000 66.2000 86.6000 66.4000 ;
	    RECT 81.2000 65.2000 82.6000 66.2000 ;
	    RECT 78.0000 62.2000 78.8000 64.2000 ;
	    RECT 81.8000 62.2000 82.6000 65.2000 ;
	    RECT 86.0000 62.2000 86.8000 66.2000 ;
	    RECT 89.2000 65.6000 90.0000 66.4000 ;
	    RECT 89.4000 64.2000 90.0000 65.6000 ;
	    RECT 92.4000 70.4000 93.0000 71.8000 ;
	    RECT 95.6000 71.6000 96.2000 75.8000 ;
	    RECT 93.8000 71.0000 96.2000 71.6000 ;
	    RECT 92.4000 69.6000 93.2000 70.4000 ;
	    RECT 92.4000 66.2000 93.0000 69.6000 ;
	    RECT 93.8000 67.6000 94.4000 71.0000 ;
	    RECT 93.6000 67.4000 94.4000 67.6000 ;
	    RECT 93.6000 67.0000 96.6000 67.4000 ;
	    RECT 93.6000 66.8000 97.8000 67.0000 ;
	    RECT 96.0000 66.4000 97.8000 66.8000 ;
	    RECT 97.2000 66.2000 97.8000 66.4000 ;
	    RECT 92.4000 65.2000 93.8000 66.2000 ;
	    RECT 93.0000 64.4000 93.8000 65.2000 ;
	    RECT 89.2000 62.2000 90.0000 64.2000 ;
	    RECT 92.4000 63.6000 93.8000 64.4000 ;
	    RECT 93.0000 62.2000 93.8000 63.6000 ;
	    RECT 97.2000 62.2000 98.0000 66.2000 ;
	    RECT 1.2000 55.6000 2.0000 57.2000 ;
	    RECT 2.8000 42.2000 3.6000 59.8000 ;
	    RECT 4.4000 54.3000 5.2000 59.8000 ;
	    RECT 6.0000 55.6000 6.8000 57.2000 ;
	    RECT 10.2000 56.4000 11.0000 59.8000 ;
	    RECT 9.2000 55.8000 11.0000 56.4000 ;
	    RECT 13.0000 56.4000 13.8000 59.8000 ;
	    RECT 19.8000 56.4000 20.6000 59.8000 ;
	    RECT 13.0000 55.8000 14.8000 56.4000 ;
	    RECT 7.6000 54.3000 8.4000 55.2000 ;
	    RECT 4.4000 53.7000 8.4000 54.3000 ;
	    RECT 4.4000 42.2000 5.2000 53.7000 ;
	    RECT 7.6000 53.6000 8.4000 53.7000 ;
	    RECT 9.2000 42.2000 10.0000 55.8000 ;
	    RECT 14.0000 52.3000 14.8000 55.8000 ;
	    RECT 18.8000 55.8000 20.6000 56.4000 ;
	    RECT 22.0000 55.8000 22.8000 59.8000 ;
	    RECT 26.2000 56.8000 27.0000 59.8000 ;
	    RECT 26.2000 55.8000 27.6000 56.8000 ;
	    RECT 33.8000 56.4000 34.6000 59.8000 ;
	    RECT 38.6000 58.4000 39.4000 59.8000 ;
	    RECT 38.0000 57.6000 39.4000 58.4000 ;
	    RECT 38.6000 56.4000 39.4000 57.6000 ;
	    RECT 33.8000 55.8000 35.6000 56.4000 ;
	    RECT 38.6000 55.8000 40.4000 56.4000 ;
	    RECT 15.6000 53.6000 16.4000 55.2000 ;
	    RECT 17.2000 53.6000 18.0000 55.2000 ;
	    RECT 10.9000 51.7000 14.8000 52.3000 ;
	    RECT 10.9000 50.4000 11.5000 51.7000 ;
	    RECT 10.8000 48.8000 11.6000 50.4000 ;
	    RECT 12.4000 48.8000 13.2000 50.4000 ;
	    RECT 14.0000 42.2000 14.8000 51.7000 ;
	    RECT 17.2000 48.3000 18.0000 48.4000 ;
	    RECT 18.8000 48.3000 19.6000 55.8000 ;
	    RECT 22.2000 55.6000 22.8000 55.8000 ;
	    RECT 22.2000 55.2000 24.0000 55.6000 ;
	    RECT 22.2000 55.0000 26.4000 55.2000 ;
	    RECT 23.4000 54.6000 26.4000 55.0000 ;
	    RECT 25.6000 54.4000 26.4000 54.6000 ;
	    RECT 20.4000 54.3000 21.2000 54.4000 ;
	    RECT 22.0000 54.3000 22.8000 54.4000 ;
	    RECT 20.4000 53.7000 22.8000 54.3000 ;
	    RECT 24.0000 53.8000 24.8000 54.0000 ;
	    RECT 20.4000 53.6000 21.2000 53.7000 ;
	    RECT 22.0000 52.8000 22.8000 53.7000 ;
	    RECT 23.8000 53.2000 24.8000 53.8000 ;
	    RECT 23.8000 52.4000 24.4000 53.2000 ;
	    RECT 23.6000 51.6000 24.4000 52.4000 ;
	    RECT 25.6000 51.0000 26.2000 54.4000 ;
	    RECT 27.0000 52.4000 27.6000 55.8000 ;
	    RECT 26.8000 51.6000 27.6000 52.4000 ;
	    RECT 23.8000 50.4000 26.2000 51.0000 ;
	    RECT 20.4000 48.8000 21.2000 50.4000 ;
	    RECT 17.2000 47.7000 19.6000 48.3000 ;
	    RECT 17.2000 47.6000 18.0000 47.7000 ;
	    RECT 18.8000 42.2000 19.6000 47.7000 ;
	    RECT 23.8000 46.2000 24.4000 50.4000 ;
	    RECT 27.0000 50.3000 27.6000 51.6000 ;
	    RECT 33.2000 50.3000 34.0000 50.4000 ;
	    RECT 26.9000 50.2000 34.0000 50.3000 ;
	    RECT 23.6000 42.2000 24.4000 46.2000 ;
	    RECT 26.8000 49.7000 34.0000 50.2000 ;
	    RECT 26.8000 42.2000 27.6000 49.7000 ;
	    RECT 33.2000 48.8000 34.0000 49.7000 ;
	    RECT 34.8000 42.2000 35.6000 55.8000 ;
	    RECT 36.4000 54.3000 37.2000 55.2000 ;
	    RECT 39.6000 54.3000 40.4000 55.8000 ;
	    RECT 36.4000 53.7000 40.4000 54.3000 ;
	    RECT 36.4000 53.6000 37.2000 53.7000 ;
	    RECT 38.0000 48.8000 38.8000 50.4000 ;
	    RECT 39.6000 42.2000 40.4000 53.7000 ;
	    RECT 41.2000 54.3000 42.0000 55.2000 ;
	    RECT 42.8000 54.3000 43.6000 59.8000 ;
	    RECT 44.4000 55.6000 45.2000 57.2000 ;
	    RECT 46.6000 56.4000 47.4000 59.8000 ;
	    RECT 46.6000 55.8000 48.4000 56.4000 ;
	    RECT 41.2000 53.7000 43.6000 54.3000 ;
	    RECT 41.2000 53.6000 42.0000 53.7000 ;
	    RECT 42.8000 42.2000 43.6000 53.7000 ;
	    RECT 44.4000 52.3000 45.2000 52.4000 ;
	    RECT 47.6000 52.3000 48.4000 55.8000 ;
	    RECT 49.2000 53.6000 50.0000 55.2000 ;
	    RECT 44.4000 51.7000 48.4000 52.3000 ;
	    RECT 44.4000 51.6000 45.2000 51.7000 ;
	    RECT 46.0000 48.8000 46.8000 50.4000 ;
	    RECT 47.6000 42.2000 48.4000 51.7000 ;
	    RECT 49.2000 50.3000 50.0000 50.4000 ;
	    RECT 50.8000 50.3000 51.6000 59.8000 ;
	    RECT 52.4000 55.6000 53.2000 57.2000 ;
	    RECT 54.6000 56.4000 55.4000 59.8000 ;
	    RECT 54.6000 55.8000 56.4000 56.4000 ;
	    RECT 52.4000 54.3000 53.2000 54.4000 ;
	    RECT 55.6000 54.3000 56.4000 55.8000 ;
	    RECT 52.4000 53.7000 56.4000 54.3000 ;
	    RECT 52.4000 53.6000 53.2000 53.7000 ;
	    RECT 49.2000 49.7000 51.6000 50.3000 ;
	    RECT 49.2000 49.6000 50.0000 49.7000 ;
	    RECT 50.8000 42.2000 51.6000 49.7000 ;
	    RECT 54.0000 48.8000 54.8000 50.4000 ;
	    RECT 55.6000 42.2000 56.4000 53.7000 ;
	    RECT 57.2000 54.3000 58.0000 55.2000 ;
	    RECT 58.8000 54.3000 59.6000 59.8000 ;
	    RECT 63.6000 57.8000 64.4000 59.8000 ;
	    RECT 60.4000 56.3000 61.2000 57.2000 ;
	    RECT 62.0000 56.3000 62.8000 56.4000 ;
	    RECT 60.4000 55.7000 62.8000 56.3000 ;
	    RECT 60.4000 55.6000 61.2000 55.7000 ;
	    RECT 62.0000 55.6000 62.8000 55.7000 ;
	    RECT 57.2000 53.7000 59.6000 54.3000 ;
	    RECT 57.2000 53.6000 58.0000 53.7000 ;
	    RECT 58.8000 42.2000 59.6000 53.7000 ;
	    RECT 63.6000 54.4000 64.2000 57.8000 ;
	    RECT 68.4000 57.6000 69.2000 59.8000 ;
	    RECT 65.2000 55.6000 66.0000 57.2000 ;
	    RECT 68.4000 54.4000 69.0000 57.6000 ;
	    RECT 70.0000 55.6000 70.8000 57.2000 ;
	    RECT 76.4000 55.8000 77.2000 59.8000 ;
	    RECT 80.6000 56.8000 81.4000 59.8000 ;
	    RECT 84.4000 57.8000 85.2000 59.8000 ;
	    RECT 80.6000 55.8000 82.0000 56.8000 ;
	    RECT 76.6000 55.6000 77.2000 55.8000 ;
	    RECT 76.6000 55.2000 78.4000 55.6000 ;
	    RECT 76.6000 55.0000 80.8000 55.2000 ;
	    RECT 77.8000 54.6000 80.8000 55.0000 ;
	    RECT 80.0000 54.4000 80.8000 54.6000 ;
	    RECT 63.6000 53.6000 64.4000 54.4000 ;
	    RECT 68.4000 53.6000 69.2000 54.4000 ;
	    RECT 70.0000 54.3000 70.8000 54.4000 ;
	    RECT 76.4000 54.3000 77.2000 54.4000 ;
	    RECT 70.0000 53.7000 77.2000 54.3000 ;
	    RECT 78.4000 53.8000 79.2000 54.0000 ;
	    RECT 70.0000 53.6000 70.8000 53.7000 ;
	    RECT 60.4000 52.3000 61.2000 52.4000 ;
	    RECT 62.0000 52.3000 62.8000 52.4000 ;
	    RECT 60.4000 51.7000 62.8000 52.3000 ;
	    RECT 60.4000 51.6000 61.2000 51.7000 ;
	    RECT 62.0000 50.8000 62.8000 51.7000 ;
	    RECT 63.6000 52.3000 64.2000 53.6000 ;
	    RECT 66.8000 52.3000 67.6000 52.4000 ;
	    RECT 63.6000 51.7000 67.6000 52.3000 ;
	    RECT 63.6000 50.2000 64.2000 51.7000 ;
	    RECT 66.8000 50.8000 67.6000 51.7000 ;
	    RECT 68.4000 50.2000 69.0000 53.6000 ;
	    RECT 76.4000 52.8000 77.2000 53.7000 ;
	    RECT 78.2000 53.2000 79.2000 53.8000 ;
	    RECT 78.2000 52.4000 78.8000 53.2000 ;
	    RECT 78.0000 51.6000 78.8000 52.4000 ;
	    RECT 80.0000 51.0000 80.6000 54.4000 ;
	    RECT 81.4000 52.4000 82.0000 55.8000 ;
	    RECT 82.8000 55.6000 83.6000 57.2000 ;
	    RECT 84.6000 54.4000 85.2000 57.8000 ;
	    RECT 87.6000 55.2000 88.4000 59.8000 ;
	    RECT 94.0000 57.8000 94.8000 59.8000 ;
	    RECT 98.8000 57.8000 99.6000 59.8000 ;
	    RECT 94.2000 56.4000 94.8000 57.8000 ;
	    RECT 94.0000 55.6000 94.8000 56.4000 ;
	    RECT 87.6000 54.6000 89.8000 55.2000 ;
	    RECT 84.4000 54.3000 85.2000 54.4000 ;
	    RECT 86.0000 54.3000 86.8000 54.4000 ;
	    RECT 84.4000 53.7000 86.8000 54.3000 ;
	    RECT 84.4000 53.6000 85.2000 53.7000 ;
	    RECT 86.0000 53.6000 86.8000 53.7000 ;
	    RECT 81.2000 52.3000 82.0000 52.4000 ;
	    RECT 82.8000 52.3000 83.6000 52.4000 ;
	    RECT 81.2000 51.7000 83.6000 52.3000 ;
	    RECT 81.2000 51.6000 82.0000 51.7000 ;
	    RECT 82.8000 51.6000 83.6000 51.7000 ;
	    RECT 78.2000 50.4000 80.6000 51.0000 ;
	    RECT 62.6000 49.4000 64.4000 50.2000 ;
	    RECT 67.4000 49.4000 69.2000 50.2000 ;
	    RECT 62.6000 42.2000 63.4000 49.4000 ;
	    RECT 67.4000 42.2000 68.2000 49.4000 ;
	    RECT 78.2000 46.2000 78.8000 50.4000 ;
	    RECT 81.4000 50.2000 82.0000 51.6000 ;
	    RECT 84.6000 50.2000 85.2000 53.6000 ;
	    RECT 86.0000 50.8000 86.8000 52.4000 ;
	    RECT 87.6000 51.6000 88.4000 53.2000 ;
	    RECT 89.2000 51.6000 89.8000 54.6000 ;
	    RECT 94.2000 54.4000 94.8000 55.6000 ;
	    RECT 99.0000 54.4000 99.6000 57.8000 ;
	    RECT 94.0000 53.6000 94.8000 54.4000 ;
	    RECT 98.8000 53.6000 99.6000 54.4000 ;
	    RECT 89.2000 50.8000 90.4000 51.6000 ;
	    RECT 89.2000 50.2000 89.8000 50.8000 ;
	    RECT 94.2000 50.2000 94.8000 53.6000 ;
	    RECT 99.0000 50.2000 99.6000 53.6000 ;
	    RECT 78.0000 42.2000 78.8000 46.2000 ;
	    RECT 81.2000 42.2000 82.0000 50.2000 ;
	    RECT 84.4000 49.4000 86.2000 50.2000 ;
	    RECT 85.4000 42.2000 86.2000 49.4000 ;
	    RECT 87.6000 49.6000 89.8000 50.2000 ;
	    RECT 87.6000 42.2000 88.4000 49.6000 ;
	    RECT 94.0000 49.4000 95.8000 50.2000 ;
	    RECT 98.8000 49.4000 100.6000 50.2000 ;
	    RECT 95.0000 42.2000 95.8000 49.4000 ;
	    RECT 99.8000 44.4000 100.6000 49.4000 ;
	    RECT 98.8000 43.6000 100.6000 44.4000 ;
	    RECT 99.8000 42.2000 100.6000 43.6000 ;
	    RECT 1.8000 32.6000 2.6000 39.8000 ;
	    RECT 7.6000 35.8000 8.4000 39.8000 ;
	    RECT 1.8000 31.8000 3.6000 32.6000 ;
	    RECT 2.8000 28.4000 3.4000 31.8000 ;
	    RECT 7.8000 31.6000 8.4000 35.8000 ;
	    RECT 10.8000 31.8000 11.6000 39.8000 ;
	    RECT 13.0000 32.6000 13.8000 39.8000 ;
	    RECT 13.0000 31.8000 14.8000 32.6000 ;
	    RECT 7.8000 31.0000 10.2000 31.6000 ;
	    RECT 2.8000 27.6000 3.6000 28.4000 ;
	    RECT 9.6000 27.6000 10.2000 31.0000 ;
	    RECT 11.0000 30.4000 11.6000 31.8000 ;
	    RECT 10.8000 30.3000 11.6000 30.4000 ;
	    RECT 12.4000 30.3000 13.2000 31.2000 ;
	    RECT 10.8000 29.7000 13.2000 30.3000 ;
	    RECT 10.8000 29.6000 11.6000 29.7000 ;
	    RECT 12.4000 29.6000 13.2000 29.7000 ;
	    RECT 2.8000 26.4000 3.4000 27.6000 ;
	    RECT 9.6000 27.4000 10.4000 27.6000 ;
	    RECT 7.4000 27.0000 10.4000 27.4000 ;
	    RECT 6.2000 26.8000 10.4000 27.0000 ;
	    RECT 6.2000 26.4000 8.0000 26.8000 ;
	    RECT 2.8000 25.6000 3.6000 26.4000 ;
	    RECT 6.2000 26.2000 6.8000 26.4000 ;
	    RECT 11.0000 26.2000 11.6000 29.6000 ;
	    RECT 2.8000 24.2000 3.4000 25.6000 ;
	    RECT 2.8000 22.2000 3.6000 24.2000 ;
	    RECT 6.0000 22.2000 6.8000 26.2000 ;
	    RECT 10.2000 25.2000 11.6000 26.2000 ;
	    RECT 14.0000 28.4000 14.6000 31.8000 ;
	    RECT 14.0000 27.6000 14.8000 28.4000 ;
	    RECT 10.2000 22.2000 11.0000 25.2000 ;
	    RECT 14.0000 24.4000 14.6000 27.6000 ;
	    RECT 15.6000 26.3000 16.4000 26.4000 ;
	    RECT 17.2000 26.3000 18.0000 26.4000 ;
	    RECT 15.6000 25.7000 18.0000 26.3000 ;
	    RECT 15.6000 24.8000 16.4000 25.7000 ;
	    RECT 17.2000 24.8000 18.0000 25.7000 ;
	    RECT 14.0000 22.2000 14.8000 24.4000 ;
	    RECT 18.8000 22.2000 19.6000 39.8000 ;
	    RECT 22.0000 28.3000 22.8000 39.8000 ;
	    RECT 23.6000 28.3000 24.4000 28.4000 ;
	    RECT 22.0000 27.7000 24.4000 28.3000 ;
	    RECT 20.4000 24.8000 21.2000 26.4000 ;
	    RECT 22.0000 22.2000 22.8000 27.7000 ;
	    RECT 23.6000 26.8000 24.4000 27.7000 ;
	    RECT 25.2000 26.2000 26.0000 39.8000 ;
	    RECT 26.8000 31.6000 27.6000 33.2000 ;
	    RECT 34.8000 28.3000 35.6000 39.8000 ;
	    RECT 36.4000 28.3000 37.2000 28.4000 ;
	    RECT 34.8000 27.7000 37.2000 28.3000 ;
	    RECT 33.2000 26.3000 34.0000 26.4000 ;
	    RECT 25.2000 25.6000 27.0000 26.2000 ;
	    RECT 26.2000 24.3000 27.0000 25.6000 ;
	    RECT 28.5000 25.7000 34.0000 26.3000 ;
	    RECT 28.5000 24.3000 29.1000 25.7000 ;
	    RECT 33.2000 24.8000 34.0000 25.7000 ;
	    RECT 26.2000 23.7000 29.1000 24.3000 ;
	    RECT 26.2000 22.2000 27.0000 23.7000 ;
	    RECT 34.8000 22.2000 35.6000 27.7000 ;
	    RECT 36.4000 26.8000 37.2000 27.7000 ;
	    RECT 38.0000 28.3000 38.8000 39.8000 ;
	    RECT 39.6000 31.6000 40.4000 33.2000 ;
	    RECT 41.2000 28.3000 42.0000 28.4000 ;
	    RECT 38.0000 27.7000 42.0000 28.3000 ;
	    RECT 38.0000 26.2000 38.8000 27.7000 ;
	    RECT 41.2000 26.8000 42.0000 27.7000 ;
	    RECT 42.8000 26.2000 43.6000 39.8000 ;
	    RECT 44.4000 32.3000 45.2000 33.2000 ;
	    RECT 46.0000 32.3000 46.8000 39.8000 ;
	    RECT 44.4000 31.7000 46.8000 32.3000 ;
	    RECT 44.4000 31.6000 45.2000 31.7000 ;
	    RECT 46.0000 30.3000 46.8000 31.7000 ;
	    RECT 49.2000 30.3000 50.0000 30.4000 ;
	    RECT 46.0000 29.7000 50.0000 30.3000 ;
	    RECT 38.0000 25.6000 39.8000 26.2000 ;
	    RECT 42.8000 25.6000 44.6000 26.2000 ;
	    RECT 39.0000 22.2000 39.8000 25.6000 ;
	    RECT 43.8000 22.2000 44.6000 25.6000 ;
	    RECT 46.0000 22.2000 46.8000 29.7000 ;
	    RECT 49.2000 29.6000 50.0000 29.7000 ;
	    RECT 49.2000 26.8000 50.0000 28.4000 ;
	    RECT 47.6000 24.8000 48.4000 26.4000 ;
	    RECT 50.8000 26.2000 51.6000 39.8000 ;
	    RECT 52.4000 32.3000 53.2000 33.2000 ;
	    RECT 54.0000 32.3000 54.8000 39.8000 ;
	    RECT 52.4000 31.8000 54.8000 32.3000 ;
	    RECT 57.2000 35.8000 58.0000 39.8000 ;
	    RECT 52.4000 31.7000 54.7000 31.8000 ;
	    RECT 52.4000 31.6000 53.2000 31.7000 ;
	    RECT 54.0000 30.4000 54.6000 31.7000 ;
	    RECT 57.2000 31.6000 57.8000 35.8000 ;
	    RECT 60.4000 31.6000 61.2000 33.2000 ;
	    RECT 55.4000 31.0000 57.8000 31.6000 ;
	    RECT 54.0000 29.6000 54.8000 30.4000 ;
	    RECT 54.0000 26.2000 54.6000 29.6000 ;
	    RECT 55.4000 27.6000 56.0000 31.0000 ;
	    RECT 57.2000 29.6000 58.0000 30.4000 ;
	    RECT 57.2000 28.8000 57.8000 29.6000 ;
	    RECT 56.8000 28.2000 57.8000 28.8000 ;
	    RECT 56.8000 28.0000 57.6000 28.2000 ;
	    RECT 58.8000 27.6000 59.6000 29.2000 ;
	    RECT 55.2000 27.4000 56.0000 27.6000 ;
	    RECT 55.2000 27.0000 58.2000 27.4000 ;
	    RECT 55.2000 26.8000 59.4000 27.0000 ;
	    RECT 57.6000 26.4000 59.4000 26.8000 ;
	    RECT 58.8000 26.2000 59.4000 26.4000 ;
	    RECT 62.0000 26.2000 62.8000 39.8000 ;
	    RECT 63.6000 28.3000 64.4000 28.4000 ;
	    RECT 65.2000 28.3000 66.0000 39.8000 ;
	    RECT 70.0000 30.3000 70.8000 39.8000 ;
	    RECT 76.4000 34.3000 77.2000 34.4000 ;
	    RECT 71.6000 33.7000 77.2000 34.3000 ;
	    RECT 71.6000 31.6000 72.4000 33.7000 ;
	    RECT 76.4000 33.6000 77.2000 33.7000 ;
	    RECT 78.0000 31.6000 78.8000 33.2000 ;
	    RECT 78.1000 30.3000 78.7000 31.6000 ;
	    RECT 70.0000 29.7000 78.7000 30.3000 ;
	    RECT 68.4000 28.3000 69.2000 28.4000 ;
	    RECT 63.6000 27.7000 66.0000 28.3000 ;
	    RECT 63.6000 26.8000 64.4000 27.7000 ;
	    RECT 50.8000 25.6000 52.6000 26.2000 ;
	    RECT 51.8000 24.4000 52.6000 25.6000 ;
	    RECT 54.0000 25.2000 55.4000 26.2000 ;
	    RECT 51.8000 23.6000 53.2000 24.4000 ;
	    RECT 51.8000 22.2000 52.6000 23.6000 ;
	    RECT 54.6000 22.2000 55.4000 25.2000 ;
	    RECT 58.8000 22.2000 59.6000 26.2000 ;
	    RECT 61.0000 25.6000 62.8000 26.2000 ;
	    RECT 61.0000 24.4000 61.8000 25.6000 ;
	    RECT 61.0000 23.6000 62.8000 24.4000 ;
	    RECT 61.0000 22.2000 61.8000 23.6000 ;
	    RECT 65.2000 22.2000 66.0000 27.7000 ;
	    RECT 66.9000 27.7000 69.2000 28.3000 ;
	    RECT 66.9000 26.4000 67.5000 27.7000 ;
	    RECT 68.4000 26.8000 69.2000 27.7000 ;
	    RECT 66.8000 24.8000 67.6000 26.4000 ;
	    RECT 70.0000 26.2000 70.8000 29.7000 ;
	    RECT 79.6000 26.2000 80.4000 39.8000 ;
	    RECT 81.2000 26.8000 82.0000 28.4000 ;
	    RECT 70.0000 25.6000 71.8000 26.2000 ;
	    RECT 71.0000 22.2000 71.8000 25.6000 ;
	    RECT 78.6000 25.6000 80.4000 26.2000 ;
	    RECT 78.6000 22.2000 79.4000 25.6000 ;
	    RECT 82.8000 22.2000 83.6000 39.8000 ;
	    RECT 84.4000 28.3000 85.2000 28.4000 ;
	    RECT 86.0000 28.3000 86.8000 39.8000 ;
	    RECT 89.8000 32.6000 90.6000 39.8000 ;
	    RECT 89.8000 31.8000 91.6000 32.6000 ;
	    RECT 94.0000 31.8000 94.8000 39.8000 ;
	    RECT 97.2000 35.8000 98.0000 39.8000 ;
	    RECT 87.6000 30.3000 88.4000 30.4000 ;
	    RECT 89.2000 30.3000 90.0000 31.2000 ;
	    RECT 87.6000 29.7000 90.0000 30.3000 ;
	    RECT 87.6000 29.6000 88.4000 29.7000 ;
	    RECT 89.2000 29.6000 90.0000 29.7000 ;
	    RECT 84.4000 27.7000 86.8000 28.3000 ;
	    RECT 84.4000 27.6000 85.2000 27.7000 ;
	    RECT 84.4000 24.8000 85.2000 26.4000 ;
	    RECT 86.0000 22.2000 86.8000 27.7000 ;
	    RECT 90.8000 28.4000 91.4000 31.8000 ;
	    RECT 94.0000 30.4000 94.6000 31.8000 ;
	    RECT 97.2000 31.6000 97.8000 35.8000 ;
	    RECT 95.4000 31.0000 97.8000 31.6000 ;
	    RECT 94.0000 29.6000 94.8000 30.4000 ;
	    RECT 90.8000 27.6000 91.6000 28.4000 ;
	    RECT 87.6000 24.8000 88.4000 26.4000 ;
	    RECT 90.8000 24.4000 91.4000 27.6000 ;
	    RECT 92.4000 24.8000 93.2000 26.4000 ;
	    RECT 94.0000 26.2000 94.6000 29.6000 ;
	    RECT 95.4000 27.6000 96.0000 31.0000 ;
	    RECT 95.2000 27.4000 96.0000 27.6000 ;
	    RECT 95.2000 27.0000 98.2000 27.4000 ;
	    RECT 95.2000 26.8000 99.4000 27.0000 ;
	    RECT 97.6000 26.4000 99.4000 26.8000 ;
	    RECT 98.8000 26.2000 99.4000 26.4000 ;
	    RECT 94.0000 25.2000 95.4000 26.2000 ;
	    RECT 90.8000 22.2000 91.6000 24.4000 ;
	    RECT 94.6000 22.2000 95.4000 25.2000 ;
	    RECT 98.8000 22.2000 99.6000 26.2000 ;
	    RECT 4.4000 15.2000 5.2000 19.8000 ;
	    RECT 7.6000 17.8000 8.4000 19.8000 ;
	    RECT 12.4000 17.8000 13.2000 19.8000 ;
	    RECT 6.0000 15.6000 6.8000 17.2000 ;
	    RECT 3.0000 14.6000 5.2000 15.2000 ;
	    RECT 3.0000 11.6000 3.6000 14.6000 ;
	    RECT 7.8000 14.4000 8.4000 17.8000 ;
	    RECT 10.8000 15.6000 11.6000 17.2000 ;
	    RECT 12.6000 16.4000 13.2000 17.8000 ;
	    RECT 12.4000 15.6000 13.2000 16.4000 ;
	    RECT 15.6000 15.8000 16.4000 19.8000 ;
	    RECT 19.8000 18.4000 20.6000 19.8000 ;
	    RECT 19.8000 17.6000 21.2000 18.4000 ;
	    RECT 19.8000 16.8000 20.6000 17.6000 ;
	    RECT 19.8000 15.8000 21.2000 16.8000 ;
	    RECT 12.6000 14.4000 13.2000 15.6000 ;
	    RECT 15.8000 15.6000 16.4000 15.8000 ;
	    RECT 15.8000 15.2000 17.6000 15.6000 ;
	    RECT 15.8000 15.0000 20.0000 15.2000 ;
	    RECT 17.0000 14.6000 20.0000 15.0000 ;
	    RECT 19.2000 14.4000 20.0000 14.6000 ;
	    RECT 7.6000 13.6000 8.4000 14.4000 ;
	    RECT 12.4000 13.6000 13.2000 14.4000 ;
	    RECT 4.4000 12.3000 5.2000 13.2000 ;
	    RECT 7.8000 12.3000 8.4000 13.6000 ;
	    RECT 4.4000 11.7000 8.4000 12.3000 ;
	    RECT 4.4000 11.6000 5.2000 11.7000 ;
	    RECT 2.4000 10.8000 3.6000 11.6000 ;
	    RECT 3.0000 10.2000 3.6000 10.8000 ;
	    RECT 7.8000 10.2000 8.4000 11.7000 ;
	    RECT 9.2000 10.8000 10.0000 12.4000 ;
	    RECT 12.6000 10.2000 13.2000 13.6000 ;
	    RECT 15.6000 12.8000 16.4000 14.4000 ;
	    RECT 17.6000 13.8000 18.4000 14.0000 ;
	    RECT 17.4000 13.2000 18.4000 13.8000 ;
	    RECT 17.4000 12.4000 18.0000 13.2000 ;
	    RECT 14.0000 10.8000 14.8000 12.4000 ;
	    RECT 17.2000 11.6000 18.0000 12.4000 ;
	    RECT 19.2000 11.0000 19.8000 14.4000 ;
	    RECT 20.6000 12.4000 21.2000 15.8000 ;
	    RECT 25.2000 15.2000 26.0000 19.8000 ;
	    RECT 33.2000 17.8000 34.0000 19.8000 ;
	    RECT 31.6000 15.6000 32.4000 17.2000 ;
	    RECT 20.4000 11.6000 21.2000 12.4000 ;
	    RECT 23.8000 14.6000 26.0000 15.2000 ;
	    RECT 23.8000 11.6000 24.4000 14.6000 ;
	    RECT 33.4000 14.4000 34.0000 17.8000 ;
	    RECT 37.0000 16.8000 37.8000 19.8000 ;
	    RECT 33.2000 13.6000 34.0000 14.4000 ;
	    RECT 25.2000 12.3000 26.0000 13.2000 ;
	    RECT 33.4000 12.3000 34.0000 13.6000 ;
	    RECT 36.4000 15.8000 37.8000 16.8000 ;
	    RECT 41.2000 15.8000 42.0000 19.8000 ;
	    RECT 44.4000 17.8000 45.2000 19.8000 ;
	    RECT 49.2000 17.8000 50.0000 19.8000 ;
	    RECT 36.4000 12.4000 37.0000 15.8000 ;
	    RECT 41.2000 15.6000 41.8000 15.8000 ;
	    RECT 40.0000 15.2000 41.8000 15.6000 ;
	    RECT 37.6000 15.0000 41.8000 15.2000 ;
	    RECT 37.6000 14.6000 40.6000 15.0000 ;
	    RECT 37.6000 14.4000 38.4000 14.6000 ;
	    RECT 44.4000 14.4000 45.0000 17.8000 ;
	    RECT 46.0000 15.6000 46.8000 17.2000 ;
	    RECT 47.6000 15.6000 48.4000 17.2000 ;
	    RECT 49.4000 14.4000 50.0000 17.8000 ;
	    RECT 54.0000 17.8000 54.8000 19.8000 ;
	    RECT 52.4000 16.3000 53.2000 16.4000 ;
	    RECT 54.0000 16.3000 54.6000 17.8000 ;
	    RECT 52.4000 15.7000 54.7000 16.3000 ;
	    RECT 57.2000 15.8000 58.0000 19.8000 ;
	    RECT 61.4000 18.4000 62.2000 19.8000 ;
	    RECT 61.4000 17.6000 62.8000 18.4000 ;
	    RECT 61.4000 16.8000 62.2000 17.6000 ;
	    RECT 61.4000 15.8000 62.8000 16.8000 ;
	    RECT 64.2000 16.4000 65.0000 19.8000 ;
	    RECT 64.2000 15.8000 66.0000 16.4000 ;
	    RECT 52.4000 15.6000 53.2000 15.7000 ;
	    RECT 25.2000 11.7000 34.0000 12.3000 ;
	    RECT 25.2000 11.6000 26.0000 11.7000 ;
	    RECT 17.4000 10.4000 19.8000 11.0000 ;
	    RECT 3.0000 9.6000 5.2000 10.2000 ;
	    RECT 4.4000 2.2000 5.2000 9.6000 ;
	    RECT 7.6000 9.4000 9.4000 10.2000 ;
	    RECT 12.4000 9.4000 14.2000 10.2000 ;
	    RECT 8.6000 2.2000 9.4000 9.4000 ;
	    RECT 13.4000 2.2000 14.2000 9.4000 ;
	    RECT 17.4000 6.2000 18.0000 10.4000 ;
	    RECT 20.6000 10.2000 21.2000 11.6000 ;
	    RECT 23.2000 10.8000 24.4000 11.6000 ;
	    RECT 17.2000 2.2000 18.0000 6.2000 ;
	    RECT 20.4000 2.2000 21.2000 10.2000 ;
	    RECT 23.8000 10.2000 24.4000 10.8000 ;
	    RECT 33.4000 10.2000 34.0000 11.7000 ;
	    RECT 34.8000 12.3000 35.6000 12.4000 ;
	    RECT 36.4000 12.3000 37.2000 12.4000 ;
	    RECT 34.8000 11.7000 37.2000 12.3000 ;
	    RECT 34.8000 10.8000 35.6000 11.7000 ;
	    RECT 36.4000 11.6000 37.2000 11.7000 ;
	    RECT 36.4000 10.2000 37.0000 11.6000 ;
	    RECT 37.8000 11.0000 38.4000 14.4000 ;
	    RECT 39.2000 13.8000 40.0000 14.0000 ;
	    RECT 39.2000 13.2000 40.2000 13.8000 ;
	    RECT 39.6000 12.4000 40.2000 13.2000 ;
	    RECT 41.2000 12.8000 42.0000 14.4000 ;
	    RECT 42.8000 14.3000 43.6000 14.4000 ;
	    RECT 44.4000 14.3000 45.2000 14.4000 ;
	    RECT 42.8000 13.7000 45.2000 14.3000 ;
	    RECT 42.8000 13.6000 43.6000 13.7000 ;
	    RECT 44.4000 13.6000 45.2000 13.7000 ;
	    RECT 49.2000 13.6000 50.0000 14.4000 ;
	    RECT 39.6000 11.6000 40.4000 12.4000 ;
	    RECT 37.8000 10.4000 40.2000 11.0000 ;
	    RECT 42.8000 10.8000 43.6000 12.4000 ;
	    RECT 23.8000 9.6000 26.0000 10.2000 ;
	    RECT 25.2000 2.2000 26.0000 9.6000 ;
	    RECT 33.2000 9.4000 35.0000 10.2000 ;
	    RECT 34.2000 2.2000 35.0000 9.4000 ;
	    RECT 36.4000 2.2000 37.2000 10.2000 ;
	    RECT 39.6000 6.2000 40.2000 10.4000 ;
	    RECT 44.4000 10.2000 45.0000 13.6000 ;
	    RECT 49.4000 12.4000 50.0000 13.6000 ;
	    RECT 54.0000 14.4000 54.6000 15.7000 ;
	    RECT 57.4000 15.6000 58.0000 15.8000 ;
	    RECT 57.4000 15.2000 59.2000 15.6000 ;
	    RECT 57.4000 15.0000 61.6000 15.2000 ;
	    RECT 58.6000 14.6000 61.6000 15.0000 ;
	    RECT 60.8000 14.4000 61.6000 14.6000 ;
	    RECT 54.0000 13.6000 54.8000 14.4000 ;
	    RECT 49.2000 11.6000 50.0000 12.4000 ;
	    RECT 49.4000 10.2000 50.0000 11.6000 ;
	    RECT 50.8000 10.8000 51.6000 12.4000 ;
	    RECT 54.0000 10.2000 54.6000 13.6000 ;
	    RECT 60.8000 11.0000 61.4000 14.4000 ;
	    RECT 62.2000 12.4000 62.8000 15.8000 ;
	    RECT 62.0000 11.6000 62.8000 12.4000 ;
	    RECT 59.0000 10.4000 61.4000 11.0000 ;
	    RECT 43.4000 9.4000 45.2000 10.2000 ;
	    RECT 49.2000 9.4000 51.0000 10.2000 ;
	    RECT 39.6000 2.2000 40.4000 6.2000 ;
	    RECT 43.4000 2.2000 44.2000 9.4000 ;
	    RECT 50.2000 2.2000 51.0000 9.4000 ;
	    RECT 53.0000 9.4000 54.8000 10.2000 ;
	    RECT 53.0000 2.2000 53.8000 9.4000 ;
	    RECT 59.0000 6.2000 59.6000 10.4000 ;
	    RECT 62.2000 10.2000 62.8000 11.6000 ;
	    RECT 65.2000 12.3000 66.0000 15.8000 ;
	    RECT 68.4000 15.2000 69.2000 19.8000 ;
	    RECT 66.8000 13.6000 67.6000 15.2000 ;
	    RECT 68.4000 14.6000 70.6000 15.2000 ;
	    RECT 68.4000 12.3000 69.2000 13.2000 ;
	    RECT 65.2000 11.7000 69.2000 12.3000 ;
	    RECT 58.8000 2.2000 59.6000 6.2000 ;
	    RECT 62.0000 2.2000 62.8000 10.2000 ;
	    RECT 63.6000 8.8000 64.4000 10.4000 ;
	    RECT 65.2000 2.2000 66.0000 11.7000 ;
	    RECT 68.4000 11.6000 69.2000 11.7000 ;
	    RECT 70.0000 11.6000 70.6000 14.6000 ;
	    RECT 73.2000 14.3000 74.0000 14.4000 ;
	    RECT 78.0000 14.3000 78.8000 19.8000 ;
	    RECT 82.8000 17.8000 83.6000 19.8000 ;
	    RECT 79.6000 15.6000 80.4000 17.2000 ;
	    RECT 81.2000 15.6000 82.0000 17.2000 ;
	    RECT 83.0000 16.3000 83.6000 17.8000 ;
	    RECT 84.4000 16.3000 85.2000 16.4000 ;
	    RECT 82.9000 15.7000 85.2000 16.3000 ;
	    RECT 86.0000 15.8000 86.8000 19.8000 ;
	    RECT 90.2000 16.8000 91.0000 19.8000 ;
	    RECT 94.0000 17.8000 94.8000 19.8000 ;
	    RECT 90.2000 15.8000 91.6000 16.8000 ;
	    RECT 83.0000 14.4000 83.6000 15.7000 ;
	    RECT 84.4000 15.6000 85.2000 15.7000 ;
	    RECT 86.2000 15.6000 86.8000 15.8000 ;
	    RECT 86.2000 15.2000 88.0000 15.6000 ;
	    RECT 86.2000 15.0000 90.4000 15.2000 ;
	    RECT 87.4000 14.6000 90.4000 15.0000 ;
	    RECT 89.6000 14.4000 90.4000 14.6000 ;
	    RECT 73.2000 13.7000 78.8000 14.3000 ;
	    RECT 73.2000 13.6000 74.0000 13.7000 ;
	    RECT 70.0000 10.8000 71.2000 11.6000 ;
	    RECT 70.0000 10.2000 70.6000 10.8000 ;
	    RECT 68.4000 9.6000 70.6000 10.2000 ;
	    RECT 68.4000 2.2000 69.2000 9.6000 ;
	    RECT 78.0000 2.2000 78.8000 13.7000 ;
	    RECT 82.8000 13.6000 83.6000 14.4000 ;
	    RECT 83.0000 10.2000 83.6000 13.6000 ;
	    RECT 86.0000 12.8000 86.8000 14.4000 ;
	    RECT 88.0000 13.8000 88.8000 14.0000 ;
	    RECT 87.8000 13.2000 88.8000 13.8000 ;
	    RECT 87.8000 12.4000 88.4000 13.2000 ;
	    RECT 84.4000 10.8000 85.2000 12.4000 ;
	    RECT 87.6000 11.6000 88.4000 12.4000 ;
	    RECT 89.6000 11.0000 90.2000 14.4000 ;
	    RECT 91.0000 12.4000 91.6000 15.8000 ;
	    RECT 94.0000 14.4000 94.6000 17.8000 ;
	    RECT 95.6000 15.6000 96.4000 17.2000 ;
	    RECT 97.2000 15.2000 98.0000 19.8000 ;
	    RECT 97.2000 14.6000 99.4000 15.2000 ;
	    RECT 94.0000 13.6000 94.8000 14.4000 ;
	    RECT 90.8000 12.3000 91.6000 12.4000 ;
	    RECT 92.4000 12.3000 93.2000 12.4000 ;
	    RECT 90.8000 11.7000 93.2000 12.3000 ;
	    RECT 90.8000 11.6000 91.6000 11.7000 ;
	    RECT 87.8000 10.4000 90.2000 11.0000 ;
	    RECT 82.8000 9.4000 84.6000 10.2000 ;
	    RECT 83.8000 2.2000 84.6000 9.4000 ;
	    RECT 87.8000 6.2000 88.4000 10.4000 ;
	    RECT 91.0000 10.2000 91.6000 11.6000 ;
	    RECT 92.4000 10.8000 93.2000 11.7000 ;
	    RECT 94.0000 12.3000 94.6000 13.6000 ;
	    RECT 97.2000 12.3000 98.0000 13.2000 ;
	    RECT 94.0000 11.7000 98.0000 12.3000 ;
	    RECT 94.0000 10.2000 94.6000 11.7000 ;
	    RECT 97.2000 11.6000 98.0000 11.7000 ;
	    RECT 98.8000 11.6000 99.4000 14.6000 ;
	    RECT 98.8000 10.8000 100.0000 11.6000 ;
	    RECT 98.8000 10.2000 99.4000 10.8000 ;
	    RECT 87.6000 2.2000 88.4000 6.2000 ;
	    RECT 90.8000 2.2000 91.6000 10.2000 ;
	    RECT 93.0000 9.4000 94.8000 10.2000 ;
	    RECT 97.2000 9.6000 99.4000 10.2000 ;
	    RECT 93.0000 2.2000 93.8000 9.4000 ;
	    RECT 97.2000 2.2000 98.0000 9.6000 ;
         LAYER metal2 ;
	    RECT 17.2000 73.6000 18.0000 74.4000 ;
	    RECT 47.6000 74.3000 48.4000 74.4000 ;
	    RECT 46.1000 73.7000 48.4000 74.3000 ;
	    RECT 12.4000 69.6000 13.2000 70.4000 ;
	    RECT 15.6000 69.6000 16.4000 70.4000 ;
	    RECT 17.3000 70.3000 17.9000 73.6000 ;
	    RECT 22.0000 71.6000 22.8000 72.4000 ;
	    RECT 33.2000 71.6000 34.0000 72.4000 ;
	    RECT 33.3000 70.4000 33.9000 71.6000 ;
	    RECT 46.1000 70.4000 46.7000 73.7000 ;
	    RECT 47.6000 73.6000 48.4000 73.7000 ;
	    RECT 55.6000 71.6000 56.4000 72.4000 ;
	    RECT 62.0000 71.6000 62.8000 72.4000 ;
	    RECT 78.0000 71.6000 78.8000 72.4000 ;
	    RECT 55.7000 70.4000 56.3000 71.6000 ;
	    RECT 62.1000 70.4000 62.7000 71.6000 ;
	    RECT 18.8000 70.3000 19.6000 70.4000 ;
	    RECT 17.3000 69.7000 19.6000 70.3000 ;
	    RECT 18.8000 69.6000 19.6000 69.7000 ;
	    RECT 23.6000 69.6000 24.4000 70.4000 ;
	    RECT 33.2000 69.6000 34.0000 70.4000 ;
	    RECT 46.0000 69.6000 46.8000 70.4000 ;
	    RECT 47.6000 69.6000 48.4000 70.4000 ;
	    RECT 50.8000 69.6000 51.6000 70.4000 ;
	    RECT 55.6000 69.6000 56.4000 70.4000 ;
	    RECT 62.0000 69.6000 62.8000 70.4000 ;
	    RECT 76.4000 69.6000 77.2000 70.4000 ;
	    RECT 81.2000 69.6000 82.0000 70.4000 ;
	    RECT 76.5000 68.4000 77.1000 69.6000 ;
	    RECT 81.3000 68.4000 81.9000 69.6000 ;
	    RECT 6.0000 67.6000 6.8000 68.4000 ;
	    RECT 17.2000 68.3000 18.0000 68.4000 ;
	    RECT 15.7000 67.7000 18.0000 68.3000 ;
	    RECT 1.2000 65.6000 2.0000 66.4000 ;
	    RECT 1.3000 64.4000 1.9000 65.6000 ;
	    RECT 1.2000 63.6000 2.0000 64.4000 ;
	    RECT 1.3000 56.4000 1.9000 63.6000 ;
	    RECT 6.1000 56.4000 6.7000 67.6000 ;
	    RECT 12.4000 65.6000 13.2000 66.4000 ;
	    RECT 12.5000 64.4000 13.1000 65.6000 ;
	    RECT 12.4000 63.6000 13.2000 64.4000 ;
	    RECT 1.2000 55.6000 2.0000 56.4000 ;
	    RECT 6.0000 55.6000 6.8000 56.4000 ;
	    RECT 6.1000 54.4000 6.7000 55.6000 ;
	    RECT 15.7000 54.4000 16.3000 67.7000 ;
	    RECT 17.2000 67.6000 18.0000 67.7000 ;
	    RECT 26.8000 67.6000 27.6000 68.4000 ;
	    RECT 38.0000 67.6000 38.8000 68.4000 ;
	    RECT 62.0000 67.6000 62.8000 68.4000 ;
	    RECT 76.4000 67.6000 77.2000 68.4000 ;
	    RECT 81.2000 67.6000 82.0000 68.4000 ;
	    RECT 26.9000 66.4000 27.5000 67.6000 ;
	    RECT 25.2000 65.6000 26.0000 66.4000 ;
	    RECT 26.8000 65.6000 27.6000 66.4000 ;
	    RECT 36.4000 65.6000 37.2000 66.4000 ;
	    RECT 38.1000 58.4000 38.7000 67.6000 ;
	    RECT 50.8000 65.6000 51.6000 66.4000 ;
	    RECT 60.4000 65.6000 61.2000 66.4000 ;
	    RECT 44.4000 63.6000 45.2000 64.4000 ;
	    RECT 60.4000 63.6000 61.2000 64.4000 ;
	    RECT 38.0000 57.6000 38.8000 58.4000 ;
	    RECT 44.5000 56.4000 45.1000 63.6000 ;
	    RECT 44.4000 55.6000 45.2000 56.4000 ;
	    RECT 52.4000 55.6000 53.2000 56.4000 ;
	    RECT 6.0000 53.6000 6.8000 54.4000 ;
	    RECT 15.6000 53.6000 16.4000 54.4000 ;
	    RECT 17.2000 53.6000 18.0000 54.4000 ;
	    RECT 20.4000 53.6000 21.2000 54.4000 ;
	    RECT 49.2000 53.6000 50.0000 54.4000 ;
	    RECT 52.4000 53.6000 53.2000 54.4000 ;
	    RECT 20.5000 50.4000 21.1000 53.6000 ;
	    RECT 60.5000 52.4000 61.1000 63.6000 ;
	    RECT 62.1000 56.4000 62.7000 67.6000 ;
	    RECT 70.0000 65.6000 70.8000 66.4000 ;
	    RECT 79.6000 65.6000 80.4000 66.4000 ;
	    RECT 89.2000 65.6000 90.0000 66.4000 ;
	    RECT 63.6000 63.6000 64.4000 64.4000 ;
	    RECT 92.4000 63.6000 93.2000 64.4000 ;
	    RECT 62.0000 55.6000 62.8000 56.4000 ;
	    RECT 23.6000 51.6000 24.4000 52.4000 ;
	    RECT 44.4000 51.6000 45.2000 52.4000 ;
	    RECT 60.4000 51.6000 61.2000 52.4000 ;
	    RECT 23.7000 50.4000 24.3000 51.6000 ;
	    RECT 44.5000 50.4000 45.1000 51.6000 ;
	    RECT 63.7000 50.4000 64.3000 63.6000 ;
	    RECT 68.4000 57.6000 69.2000 58.4000 ;
	    RECT 82.8000 57.6000 83.6000 58.4000 ;
	    RECT 82.9000 56.4000 83.5000 57.6000 ;
	    RECT 65.2000 55.6000 66.0000 56.4000 ;
	    RECT 70.0000 55.6000 70.8000 56.4000 ;
	    RECT 82.8000 55.6000 83.6000 56.4000 ;
	    RECT 94.0000 55.6000 94.8000 56.4000 ;
	    RECT 70.1000 54.4000 70.7000 55.6000 ;
	    RECT 70.0000 53.6000 70.8000 54.4000 ;
	    RECT 86.0000 54.3000 86.8000 54.4000 ;
	    RECT 86.0000 53.7000 88.3000 54.3000 ;
	    RECT 86.0000 53.6000 86.8000 53.7000 ;
	    RECT 87.7000 52.4000 88.3000 53.7000 ;
	    RECT 66.8000 51.6000 67.6000 52.4000 ;
	    RECT 78.0000 51.6000 78.8000 52.4000 ;
	    RECT 82.8000 51.6000 83.6000 52.4000 ;
	    RECT 86.0000 51.6000 86.8000 52.4000 ;
	    RECT 87.6000 51.6000 88.4000 52.4000 ;
	    RECT 2.8000 49.6000 3.6000 50.4000 ;
	    RECT 12.4000 49.6000 13.2000 50.4000 ;
	    RECT 20.4000 50.3000 21.2000 50.4000 ;
	    RECT 18.9000 49.7000 21.2000 50.3000 ;
	    RECT 17.2000 47.6000 18.0000 48.4000 ;
	    RECT 9.2000 43.6000 10.0000 44.4000 ;
	    RECT 2.8000 25.6000 3.6000 26.4000 ;
	    RECT 6.0000 15.6000 6.8000 16.4000 ;
	    RECT 9.3000 16.3000 9.9000 43.6000 ;
	    RECT 17.3000 32.4000 17.9000 47.6000 ;
	    RECT 18.9000 38.4000 19.5000 49.7000 ;
	    RECT 20.4000 49.6000 21.2000 49.7000 ;
	    RECT 23.6000 49.6000 24.4000 50.4000 ;
	    RECT 38.0000 49.6000 38.8000 50.4000 ;
	    RECT 44.4000 49.6000 45.2000 50.4000 ;
	    RECT 46.0000 49.6000 46.8000 50.4000 ;
	    RECT 49.2000 49.6000 50.0000 50.4000 ;
	    RECT 54.0000 49.6000 54.8000 50.4000 ;
	    RECT 63.6000 49.6000 64.4000 50.4000 ;
	    RECT 34.8000 43.6000 35.6000 44.4000 ;
	    RECT 98.8000 43.6000 99.6000 44.4000 ;
	    RECT 18.8000 37.6000 19.6000 38.4000 ;
	    RECT 34.9000 32.4000 35.5000 43.6000 ;
	    RECT 58.8000 33.6000 59.6000 34.4000 ;
	    RECT 76.4000 33.6000 77.2000 34.4000 ;
	    RECT 82.8000 33.6000 83.6000 34.4000 ;
	    RECT 17.2000 31.6000 18.0000 32.4000 ;
	    RECT 26.8000 31.6000 27.6000 32.4000 ;
	    RECT 34.8000 31.6000 35.6000 32.4000 ;
	    RECT 39.6000 31.6000 40.4000 32.4000 ;
	    RECT 42.8000 31.6000 43.6000 32.4000 ;
	    RECT 12.4000 29.6000 13.2000 30.4000 ;
	    RECT 49.2000 29.6000 50.0000 30.4000 ;
	    RECT 57.2000 29.6000 58.0000 30.4000 ;
	    RECT 12.5000 28.4000 13.1000 29.6000 ;
	    RECT 58.9000 28.4000 59.5000 33.6000 ;
	    RECT 60.4000 31.6000 61.2000 32.4000 ;
	    RECT 87.6000 29.6000 88.4000 30.4000 ;
	    RECT 94.0000 29.6000 94.8000 30.4000 ;
	    RECT 12.4000 27.6000 13.2000 28.4000 ;
	    RECT 20.4000 27.6000 21.2000 28.4000 ;
	    RECT 41.2000 27.6000 42.0000 28.4000 ;
	    RECT 49.2000 27.6000 50.0000 28.4000 ;
	    RECT 58.8000 27.6000 59.6000 28.4000 ;
	    RECT 81.2000 27.6000 82.0000 28.4000 ;
	    RECT 84.4000 27.6000 85.2000 28.4000 ;
	    RECT 20.5000 26.4000 21.1000 27.6000 ;
	    RECT 15.6000 25.6000 16.4000 26.4000 ;
	    RECT 20.4000 25.6000 21.2000 26.4000 ;
	    RECT 14.0000 23.6000 14.8000 24.4000 ;
	    RECT 10.8000 16.3000 11.6000 16.4000 ;
	    RECT 9.3000 15.7000 11.6000 16.3000 ;
	    RECT 10.8000 15.6000 11.6000 15.7000 ;
	    RECT 12.4000 15.6000 13.2000 16.4000 ;
	    RECT 10.9000 14.4000 11.5000 15.6000 ;
	    RECT 10.8000 13.6000 11.6000 14.4000 ;
	    RECT 14.1000 12.4000 14.7000 23.6000 ;
	    RECT 20.4000 17.6000 21.2000 18.4000 ;
	    RECT 41.3000 16.4000 41.9000 27.6000 ;
	    RECT 87.7000 26.4000 88.3000 29.6000 ;
	    RECT 98.9000 26.4000 99.5000 43.6000 ;
	    RECT 47.6000 25.6000 48.4000 26.4000 ;
	    RECT 66.8000 25.6000 67.6000 26.4000 ;
	    RECT 79.6000 25.6000 80.4000 26.4000 ;
	    RECT 84.4000 25.6000 85.2000 26.4000 ;
	    RECT 87.6000 25.6000 88.4000 26.4000 ;
	    RECT 92.4000 25.6000 93.2000 26.4000 ;
	    RECT 98.8000 25.6000 99.6000 26.4000 ;
	    RECT 47.7000 16.4000 48.3000 25.6000 ;
	    RECT 52.4000 23.6000 53.2000 24.4000 ;
	    RECT 62.0000 23.6000 62.8000 24.4000 ;
	    RECT 52.5000 20.4000 53.1000 23.6000 ;
	    RECT 52.4000 19.6000 53.2000 20.4000 ;
	    RECT 63.6000 19.6000 64.4000 20.4000 ;
	    RECT 50.8000 17.6000 51.6000 18.4000 ;
	    RECT 62.0000 17.6000 62.8000 18.4000 ;
	    RECT 31.6000 15.6000 32.4000 16.4000 ;
	    RECT 41.2000 15.6000 42.0000 16.4000 ;
	    RECT 46.0000 15.6000 46.8000 16.4000 ;
	    RECT 47.6000 15.6000 48.4000 16.4000 ;
	    RECT 31.7000 14.4000 32.3000 15.6000 ;
	    RECT 41.3000 14.4000 41.9000 15.6000 ;
	    RECT 15.6000 13.6000 16.4000 14.4000 ;
	    RECT 31.6000 13.6000 32.4000 14.4000 ;
	    RECT 41.2000 13.6000 42.0000 14.4000 ;
	    RECT 42.8000 13.6000 43.6000 14.4000 ;
	    RECT 50.9000 12.4000 51.5000 17.6000 ;
	    RECT 52.4000 15.6000 53.2000 16.4000 ;
	    RECT 9.2000 11.6000 10.0000 12.4000 ;
	    RECT 14.0000 11.6000 14.8000 12.4000 ;
	    RECT 17.2000 11.6000 18.0000 12.4000 ;
	    RECT 39.6000 11.6000 40.4000 12.4000 ;
	    RECT 42.8000 11.6000 43.6000 12.4000 ;
	    RECT 49.2000 11.6000 50.0000 12.4000 ;
	    RECT 50.8000 11.6000 51.6000 12.4000 ;
	    RECT 63.7000 10.4000 64.3000 19.6000 ;
	    RECT 66.9000 18.4000 67.5000 25.6000 ;
	    RECT 66.8000 17.6000 67.6000 18.4000 ;
	    RECT 79.7000 16.4000 80.3000 25.6000 ;
	    RECT 81.2000 23.6000 82.0000 24.4000 ;
	    RECT 86.0000 23.6000 86.8000 24.4000 ;
	    RECT 90.8000 23.6000 91.6000 24.4000 ;
	    RECT 81.3000 16.4000 81.9000 23.6000 ;
	    RECT 79.6000 15.6000 80.4000 16.4000 ;
	    RECT 81.2000 15.6000 82.0000 16.4000 ;
	    RECT 84.4000 15.6000 85.2000 16.4000 ;
	    RECT 86.1000 14.4000 86.7000 23.6000 ;
	    RECT 66.8000 13.6000 67.6000 14.4000 ;
	    RECT 73.2000 13.6000 74.0000 14.4000 ;
	    RECT 86.0000 13.6000 86.8000 14.4000 ;
	    RECT 90.9000 12.4000 91.5000 23.6000 ;
	    RECT 95.6000 15.6000 96.4000 16.4000 ;
	    RECT 84.4000 11.6000 85.2000 12.4000 ;
	    RECT 87.6000 11.6000 88.4000 12.4000 ;
	    RECT 90.8000 11.6000 91.6000 12.4000 ;
	    RECT 63.6000 9.6000 64.4000 10.4000 ;
         LAYER M3 ;
	    RECT 22.0000 72.3000 22.8000 72.4000 ;
	    RECT 33.2000 72.3000 34.0000 72.4000 ;
	    RECT 22.0000 71.7000 34.0000 72.3000 ;
	    RECT 22.0000 71.6000 22.8000 71.7000 ;
	    RECT 33.2000 71.6000 34.0000 71.7000 ;
	    RECT 55.6000 72.3000 56.4000 72.4000 ;
	    RECT 62.0000 72.3000 62.8000 72.4000 ;
	    RECT 78.0000 72.3000 78.8000 72.4000 ;
	    RECT 55.6000 71.7000 78.8000 72.3000 ;
	    RECT 55.6000 71.6000 56.4000 71.7000 ;
	    RECT 62.0000 71.6000 62.8000 71.7000 ;
	    RECT 78.0000 71.6000 78.8000 71.7000 ;
	    RECT 12.4000 70.3000 13.2000 70.4000 ;
	    RECT 15.6000 70.3000 16.4000 70.4000 ;
	    RECT 12.4000 69.7000 16.4000 70.3000 ;
	    RECT 12.4000 69.6000 13.2000 69.7000 ;
	    RECT 15.6000 69.6000 16.4000 69.7000 ;
	    RECT 18.8000 70.3000 19.6000 70.4000 ;
	    RECT 23.6000 70.3000 24.4000 70.4000 ;
	    RECT 18.8000 69.7000 24.4000 70.3000 ;
	    RECT 18.8000 69.6000 19.6000 69.7000 ;
	    RECT 23.6000 69.6000 24.4000 69.7000 ;
	    RECT 47.6000 70.3000 48.4000 70.4000 ;
	    RECT 50.8000 70.3000 51.6000 70.4000 ;
	    RECT 47.6000 69.7000 51.6000 70.3000 ;
	    RECT 47.6000 69.6000 48.4000 69.7000 ;
	    RECT 50.8000 69.6000 51.6000 69.7000 ;
	    RECT 6.0000 68.3000 6.8000 68.4000 ;
	    RECT 12.5000 68.3000 13.1000 69.6000 ;
	    RECT 6.0000 67.7000 13.1000 68.3000 ;
	    RECT 17.2000 68.3000 18.0000 68.4000 ;
	    RECT 26.8000 68.3000 27.6000 68.4000 ;
	    RECT 38.0000 68.3000 38.8000 68.4000 ;
	    RECT 17.2000 67.7000 38.8000 68.3000 ;
	    RECT 6.0000 67.6000 6.8000 67.7000 ;
	    RECT 17.2000 67.6000 18.0000 67.7000 ;
	    RECT 26.8000 67.6000 27.6000 67.7000 ;
	    RECT 38.0000 67.6000 38.8000 67.7000 ;
	    RECT 62.0000 68.3000 62.8000 68.4000 ;
	    RECT 76.4000 68.3000 77.2000 68.4000 ;
	    RECT 81.2000 68.3000 82.0000 68.4000 ;
	    RECT 62.0000 67.7000 82.0000 68.3000 ;
	    RECT 62.0000 67.6000 62.8000 67.7000 ;
	    RECT 76.4000 67.6000 77.2000 67.7000 ;
	    RECT 81.2000 67.6000 82.0000 67.7000 ;
	    RECT 25.2000 66.3000 26.0000 66.4000 ;
	    RECT 36.4000 66.3000 37.2000 66.4000 ;
	    RECT 25.2000 65.7000 37.2000 66.3000 ;
	    RECT 25.2000 65.6000 26.0000 65.7000 ;
	    RECT 36.4000 65.6000 37.2000 65.7000 ;
	    RECT 50.8000 66.3000 51.6000 66.4000 ;
	    RECT 60.4000 66.3000 61.2000 66.4000 ;
	    RECT 50.8000 65.7000 61.2000 66.3000 ;
	    RECT 50.8000 65.6000 51.6000 65.7000 ;
	    RECT 60.4000 65.6000 61.2000 65.7000 ;
	    RECT 70.0000 66.3000 70.8000 66.4000 ;
	    RECT 79.6000 66.3000 80.4000 66.4000 ;
	    RECT 89.2000 66.3000 90.0000 66.4000 ;
	    RECT 70.0000 65.7000 90.0000 66.3000 ;
	    RECT 70.0000 65.6000 70.8000 65.7000 ;
	    RECT 79.6000 65.6000 80.4000 65.7000 ;
	    RECT 89.2000 65.6000 90.0000 65.7000 ;
	    RECT 1.2000 64.3000 2.0000 64.4000 ;
	    RECT 12.4000 64.3000 13.2000 64.4000 ;
	    RECT 1.2000 63.7000 13.2000 64.3000 ;
	    RECT 1.2000 63.6000 2.0000 63.7000 ;
	    RECT 12.4000 63.6000 13.2000 63.7000 ;
	    RECT 44.4000 64.3000 45.2000 64.4000 ;
	    RECT 60.4000 64.3000 61.2000 64.4000 ;
	    RECT 92.4000 64.3000 93.2000 64.4000 ;
	    RECT 44.4000 63.7000 93.2000 64.3000 ;
	    RECT 44.4000 63.6000 45.2000 63.7000 ;
	    RECT 60.4000 63.6000 61.2000 63.7000 ;
	    RECT 92.4000 63.6000 93.2000 63.7000 ;
	    RECT 68.4000 58.3000 69.2000 58.4000 ;
	    RECT 82.8000 58.3000 83.6000 58.4000 ;
	    RECT 68.4000 57.7000 83.6000 58.3000 ;
	    RECT 68.4000 57.6000 69.2000 57.7000 ;
	    RECT 82.8000 57.6000 83.6000 57.7000 ;
	    RECT 52.4000 56.3000 53.2000 56.4000 ;
	    RECT 65.2000 56.3000 66.0000 56.4000 ;
	    RECT 94.0000 56.3000 94.8000 56.4000 ;
	    RECT 52.4000 55.7000 94.8000 56.3000 ;
	    RECT 52.4000 55.6000 53.2000 55.7000 ;
	    RECT 65.2000 55.6000 66.0000 55.7000 ;
	    RECT 94.0000 55.6000 94.8000 55.7000 ;
	    RECT 6.0000 54.3000 6.8000 54.4000 ;
	    RECT 17.2000 54.3000 18.0000 54.4000 ;
	    RECT 6.0000 53.7000 18.0000 54.3000 ;
	    RECT 6.0000 53.6000 6.8000 53.7000 ;
	    RECT 17.2000 53.6000 18.0000 53.7000 ;
	    RECT 49.2000 54.3000 50.0000 54.4000 ;
	    RECT 52.4000 54.3000 53.2000 54.4000 ;
	    RECT 70.0000 54.3000 70.8000 54.4000 ;
	    RECT 49.2000 53.7000 70.8000 54.3000 ;
	    RECT 49.2000 53.6000 50.0000 53.7000 ;
	    RECT 52.4000 53.6000 53.2000 53.7000 ;
	    RECT 70.0000 53.6000 70.8000 53.7000 ;
	    RECT 66.8000 52.3000 67.6000 52.4000 ;
	    RECT 78.0000 52.3000 78.8000 52.4000 ;
	    RECT 66.8000 51.7000 78.8000 52.3000 ;
	    RECT 66.8000 51.6000 67.6000 51.7000 ;
	    RECT 78.0000 51.6000 78.8000 51.7000 ;
	    RECT 82.8000 52.3000 83.6000 52.4000 ;
	    RECT 86.0000 52.3000 86.8000 52.4000 ;
	    RECT 82.8000 51.7000 86.8000 52.3000 ;
	    RECT 82.8000 51.6000 83.6000 51.7000 ;
	    RECT 86.0000 51.6000 86.8000 51.7000 ;
	    RECT 2.8000 50.3000 3.6000 50.4000 ;
	    RECT 12.4000 50.3000 13.2000 50.4000 ;
	    RECT 23.6000 50.3000 24.4000 50.4000 ;
	    RECT 2.8000 49.7000 24.4000 50.3000 ;
	    RECT 2.8000 49.6000 3.6000 49.7000 ;
	    RECT 12.4000 49.6000 13.2000 49.7000 ;
	    RECT 23.6000 49.6000 24.4000 49.7000 ;
	    RECT 38.0000 50.3000 38.8000 50.4000 ;
	    RECT 44.4000 50.3000 45.2000 50.4000 ;
	    RECT 38.0000 49.7000 45.2000 50.3000 ;
	    RECT 38.0000 49.6000 38.8000 49.7000 ;
	    RECT 44.4000 49.6000 45.2000 49.7000 ;
	    RECT 46.0000 50.3000 46.8000 50.4000 ;
	    RECT 49.2000 50.3000 50.0000 50.4000 ;
	    RECT 46.0000 49.7000 50.0000 50.3000 ;
	    RECT 46.0000 49.6000 46.8000 49.7000 ;
	    RECT 49.2000 49.6000 50.0000 49.7000 ;
	    RECT 54.0000 50.3000 54.8000 50.4000 ;
	    RECT 63.6000 50.3000 64.4000 50.4000 ;
	    RECT 54.0000 49.7000 64.4000 50.3000 ;
	    RECT 54.0000 49.6000 54.8000 49.7000 ;
	    RECT 63.6000 49.6000 64.4000 49.7000 ;
	    RECT 58.8000 34.3000 59.6000 34.4000 ;
	    RECT 76.4000 34.3000 77.2000 34.4000 ;
	    RECT 82.8000 34.3000 83.6000 34.4000 ;
	    RECT 58.8000 33.7000 83.6000 34.3000 ;
	    RECT 58.8000 33.6000 59.6000 33.7000 ;
	    RECT 76.4000 33.6000 77.2000 33.7000 ;
	    RECT 82.8000 33.6000 83.6000 33.7000 ;
	    RECT 17.2000 32.3000 18.0000 32.4000 ;
	    RECT 26.8000 32.3000 27.6000 32.4000 ;
	    RECT 17.2000 31.7000 27.6000 32.3000 ;
	    RECT 17.2000 31.6000 18.0000 31.7000 ;
	    RECT 26.8000 31.6000 27.6000 31.7000 ;
	    RECT 34.8000 32.3000 35.6000 32.4000 ;
	    RECT 39.6000 32.3000 40.4000 32.4000 ;
	    RECT 34.8000 31.7000 40.4000 32.3000 ;
	    RECT 34.8000 31.6000 35.6000 31.7000 ;
	    RECT 39.6000 31.6000 40.4000 31.7000 ;
	    RECT 42.8000 32.3000 43.6000 32.4000 ;
	    RECT 60.4000 32.3000 61.2000 32.4000 ;
	    RECT 42.8000 31.7000 61.2000 32.3000 ;
	    RECT 42.8000 31.6000 43.6000 31.7000 ;
	    RECT 60.4000 31.6000 61.2000 31.7000 ;
	    RECT 49.2000 30.3000 50.0000 30.4000 ;
	    RECT 57.2000 30.3000 58.0000 30.4000 ;
	    RECT 49.2000 29.7000 58.0000 30.3000 ;
	    RECT 49.2000 29.6000 50.0000 29.7000 ;
	    RECT 57.2000 29.6000 58.0000 29.7000 ;
	    RECT 87.6000 30.3000 88.4000 30.4000 ;
	    RECT 94.0000 30.3000 94.8000 30.4000 ;
	    RECT 87.6000 29.7000 94.8000 30.3000 ;
	    RECT 87.6000 29.6000 88.4000 29.7000 ;
	    RECT 94.0000 29.6000 94.8000 29.7000 ;
	    RECT 12.4000 28.3000 13.2000 28.4000 ;
	    RECT 20.4000 28.3000 21.2000 28.4000 ;
	    RECT 12.4000 27.7000 21.2000 28.3000 ;
	    RECT 12.4000 27.6000 13.2000 27.7000 ;
	    RECT 20.4000 27.6000 21.2000 27.7000 ;
	    RECT 41.2000 28.3000 42.0000 28.4000 ;
	    RECT 49.2000 28.3000 50.0000 28.4000 ;
	    RECT 41.2000 27.7000 50.0000 28.3000 ;
	    RECT 41.2000 27.6000 42.0000 27.7000 ;
	    RECT 49.2000 27.6000 50.0000 27.7000 ;
	    RECT 81.2000 28.3000 82.0000 28.4000 ;
	    RECT 84.4000 28.3000 85.2000 28.4000 ;
	    RECT 81.2000 27.7000 85.2000 28.3000 ;
	    RECT 81.2000 27.6000 82.0000 27.7000 ;
	    RECT 84.4000 27.6000 85.2000 27.7000 ;
	    RECT 2.8000 26.3000 3.6000 26.4000 ;
	    RECT 15.6000 26.3000 16.4000 26.4000 ;
	    RECT 2.8000 25.7000 16.4000 26.3000 ;
	    RECT 2.8000 25.6000 3.6000 25.7000 ;
	    RECT 15.6000 25.6000 16.4000 25.7000 ;
	    RECT 84.4000 26.3000 85.2000 26.4000 ;
	    RECT 92.4000 26.3000 93.2000 26.4000 ;
	    RECT 98.8000 26.3000 99.6000 26.4000 ;
	    RECT 84.4000 25.7000 99.6000 26.3000 ;
	    RECT 84.4000 25.6000 85.2000 25.7000 ;
	    RECT 92.4000 25.6000 93.2000 25.7000 ;
	    RECT 98.8000 25.6000 99.6000 25.7000 ;
	    RECT 62.0000 24.3000 62.8000 24.4000 ;
	    RECT 81.2000 24.3000 82.0000 24.4000 ;
	    RECT 86.0000 24.3000 86.8000 24.4000 ;
	    RECT 62.0000 23.7000 86.8000 24.3000 ;
	    RECT 62.0000 23.6000 62.8000 23.7000 ;
	    RECT 81.2000 23.6000 82.0000 23.7000 ;
	    RECT 86.0000 23.6000 86.8000 23.7000 ;
	    RECT 52.4000 20.3000 53.2000 20.4000 ;
	    RECT 63.6000 20.3000 64.4000 20.4000 ;
	    RECT 52.4000 19.7000 64.4000 20.3000 ;
	    RECT 52.4000 19.6000 53.2000 19.7000 ;
	    RECT 63.6000 19.6000 64.4000 19.7000 ;
	    RECT 10.8000 18.3000 11.6000 18.4000 ;
	    RECT 20.4000 18.3000 21.2000 18.4000 ;
	    RECT 10.8000 17.7000 21.2000 18.3000 ;
	    RECT 10.8000 17.6000 11.6000 17.7000 ;
	    RECT 20.4000 17.6000 21.2000 17.7000 ;
	    RECT 50.8000 18.3000 51.6000 18.4000 ;
	    RECT 62.0000 18.3000 62.8000 18.4000 ;
	    RECT 66.8000 18.3000 67.6000 18.4000 ;
	    RECT 50.8000 17.7000 67.6000 18.3000 ;
	    RECT 50.8000 17.6000 51.6000 17.7000 ;
	    RECT 62.0000 17.6000 62.8000 17.7000 ;
	    RECT 66.8000 17.6000 67.6000 17.7000 ;
	    RECT 6.0000 16.3000 6.8000 16.4000 ;
	    RECT 12.4000 16.3000 13.2000 16.4000 ;
	    RECT 6.0000 15.7000 13.2000 16.3000 ;
	    RECT 6.0000 15.6000 6.8000 15.7000 ;
	    RECT 12.4000 15.6000 13.2000 15.7000 ;
	    RECT 41.2000 16.3000 42.0000 16.4000 ;
	    RECT 46.0000 16.3000 46.8000 16.4000 ;
	    RECT 41.2000 15.7000 46.8000 16.3000 ;
	    RECT 41.2000 15.6000 42.0000 15.7000 ;
	    RECT 46.0000 15.6000 46.8000 15.7000 ;
	    RECT 47.6000 16.3000 48.4000 16.4000 ;
	    RECT 52.4000 16.3000 53.2000 16.4000 ;
	    RECT 47.6000 15.7000 53.2000 16.3000 ;
	    RECT 47.6000 15.6000 48.4000 15.7000 ;
	    RECT 52.4000 15.6000 53.2000 15.7000 ;
	    RECT 84.4000 16.3000 85.2000 16.4000 ;
	    RECT 95.6000 16.3000 96.4000 16.4000 ;
	    RECT 84.4000 15.7000 96.4000 16.3000 ;
	    RECT 84.4000 15.6000 85.2000 15.7000 ;
	    RECT 95.6000 15.6000 96.4000 15.7000 ;
	    RECT 10.8000 14.3000 11.6000 14.4000 ;
	    RECT 15.6000 14.3000 16.4000 14.4000 ;
	    RECT 10.8000 13.7000 16.4000 14.3000 ;
	    RECT 10.8000 13.6000 11.6000 13.7000 ;
	    RECT 15.6000 13.6000 16.4000 13.7000 ;
	    RECT 31.6000 14.3000 32.4000 14.4000 ;
	    RECT 42.8000 14.3000 43.6000 14.4000 ;
	    RECT 31.6000 13.7000 43.6000 14.3000 ;
	    RECT 31.6000 13.6000 32.4000 13.7000 ;
	    RECT 42.8000 13.6000 43.6000 13.7000 ;
	    RECT 66.8000 14.3000 67.6000 14.4000 ;
	    RECT 73.2000 14.3000 74.0000 14.4000 ;
	    RECT 66.8000 13.7000 74.0000 14.3000 ;
	    RECT 66.8000 13.6000 67.6000 13.7000 ;
	    RECT 73.2000 13.6000 74.0000 13.7000 ;
	    RECT 9.2000 12.3000 10.0000 12.4000 ;
	    RECT 10.8000 12.3000 11.6000 12.4000 ;
	    RECT 9.2000 11.7000 11.6000 12.3000 ;
	    RECT 9.2000 11.6000 10.0000 11.7000 ;
	    RECT 10.8000 11.6000 11.6000 11.7000 ;
	    RECT 14.0000 12.3000 14.8000 12.4000 ;
	    RECT 17.2000 12.3000 18.0000 12.4000 ;
	    RECT 14.0000 11.7000 18.0000 12.3000 ;
	    RECT 14.0000 11.6000 14.8000 11.7000 ;
	    RECT 17.2000 11.6000 18.0000 11.7000 ;
	    RECT 39.6000 12.3000 40.4000 12.4000 ;
	    RECT 42.8000 12.3000 43.6000 12.4000 ;
	    RECT 49.2000 12.3000 50.0000 12.4000 ;
	    RECT 39.6000 11.7000 50.0000 12.3000 ;
	    RECT 39.6000 11.6000 40.4000 11.7000 ;
	    RECT 42.8000 11.6000 43.6000 11.7000 ;
	    RECT 49.2000 11.6000 50.0000 11.7000 ;
	    RECT 84.4000 12.3000 85.2000 12.4000 ;
	    RECT 87.6000 12.3000 88.4000 12.4000 ;
	    RECT 90.8000 12.3000 91.6000 12.4000 ;
	    RECT 84.4000 11.7000 91.6000 12.3000 ;
	    RECT 84.4000 11.6000 85.2000 11.7000 ;
	    RECT 87.6000 11.6000 88.4000 11.7000 ;
	    RECT 90.8000 11.6000 91.6000 11.7000 ;
         LAYER M4 ;
	    RECT 10.6000 11.4000 11.8000 18.6000 ;
   END
END PPA_adder
