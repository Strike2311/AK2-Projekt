* NGSPICE file created from PPA_adder.ext - technology: scmos

.global vdd gnd 

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

.subckt PPA_adder vdd gnd sum_comp_1[0] sum_comp_1[1] sum_comp_1[2] sum_comp_1[3]
+ sum_comp_1[4] sum_comp_1[5] sum_comp_2[0] sum_comp_2[1] sum_comp_2[2] sum_comp_2[3]
+ sum_comp_2[4] sum_comp_2[5] c_in result[0] result[1] result[2] result[3] result[4]
+ result[5] c_out
XFILL_0_0_2 gnd vdd FILL
XFILL_1_1_0 gnd vdd FILL
XBUFX2_3 BUFX2_3/A gnd result[3] vdd BUFX2
XNAND2X1_13 AND2X2_4/A AND2X2_14/Y gnd NAND2X1_14/B vdd NAND2X1
XNAND2X1_2 INVX1_1/Y NAND2X1_1/Y gnd AND2X2_7/A vdd NAND2X1
XFILL_1_1_1 gnd vdd FILL
XNAND2X1_14 INVX1_13/Y NAND2X1_14/B gnd AND2X2_6/A vdd NAND2X1
XBUFX2_4 BUFX2_4/A gnd result[4] vdd BUFX2
XNAND2X1_3 AND2X2_6/A AND2X2_1/Y gnd NAND2X1_4/B vdd NAND2X1
XFILL_1_1_2 gnd vdd FILL
XBUFX2_5 BUFX2_5/A gnd result[5] vdd BUFX2
XNAND2X1_15 INVX1_12/A INVX1_8/Y gnd NAND2X1_16/B vdd NAND2X1
XNAND2X1_4 INVX1_2/Y NAND2X1_4/B gnd BUFX2_6/A vdd NAND2X1
XNAND2X1_16 INVX1_14/Y NAND2X1_16/B gnd INVX1_13/A vdd NAND2X1
XBUFX2_6 BUFX2_6/A gnd c_out vdd BUFX2
XNAND2X1_5 INVX1_1/A AND2X2_1/A gnd NAND2X1_5/Y vdd NAND2X1
XBUFX2_7 BUFX2_7/A gnd result[0] vdd BUFX2
XNAND2X1_6 INVX1_3/Y NAND2X1_5/Y gnd INVX1_2/A vdd NAND2X1
XFILL_4_1 gnd vdd FILL
XNOR2X1_1 c_in AND2X2_2/B gnd NOR2X1_2/A vdd NOR2X1
XNAND2X1_7 INVX1_5/Y c_in gnd NAND2X1_8/B vdd NAND2X1
XFILL_4_2 gnd vdd FILL
XNOR2X1_2 NOR2X1_2/A NOR2X1_2/B gnd BUFX2_7/A vdd NOR2X1
XNAND2X1_8 INVX1_4/Y NAND2X1_8/B gnd NOR2X1_3/A vdd NAND2X1
XNAND2X1_9 NOR2X1_3/A INVX1_6/Y gnd NAND2X1_9/Y vdd NAND2X1
XNOR2X1_3 NOR2X1_3/A NOR2X1_3/B gnd NOR2X1_3/Y vdd NOR2X1
XNOR2X1_4 NOR2X1_3/Y AND2X2_3/Y gnd BUFX2_1/A vdd NOR2X1
XFILL_1_0_0 gnd vdd FILL
XINVX1_10 INVX1_10/A gnd AND2X2_1/A vdd INVX1
XFILL_1_0_1 gnd vdd FILL
XNOR2X1_5 AND2X2_4/A AND2X2_4/B gnd NOR2X1_5/Y vdd NOR2X1
XINVX1_11 INVX1_11/A gnd INVX1_11/Y vdd INVX1
XNOR2X1_6 NOR2X1_5/Y AND2X2_4/Y gnd BUFX2_2/A vdd NOR2X1
XFILL_2_1_0 gnd vdd FILL
XFILL_1_0_2 gnd vdd FILL
XINVX1_12 INVX1_12/A gnd INVX1_12/Y vdd INVX1
XFILL_2_1_1 gnd vdd FILL
XINVX1_1 INVX1_1/A gnd INVX1_1/Y vdd INVX1
XNOR2X1_7 NOR2X1_7/A NOR2X1_7/B gnd NOR2X1_8/A vdd NOR2X1
XINVX1_13 INVX1_13/A gnd INVX1_13/Y vdd INVX1
XNOR2X1_8 NOR2X1_8/A NOR2X1_8/B gnd BUFX2_3/A vdd NOR2X1
XINVX1_2 INVX1_2/A gnd INVX1_2/Y vdd INVX1
XFILL_2_1_2 gnd vdd FILL
XINVX1_14 INVX1_14/A gnd INVX1_14/Y vdd INVX1
XINVX1_3 INVX1_3/A gnd INVX1_3/Y vdd INVX1
XNOR2X1_9 AND2X2_6/A AND2X2_6/B gnd NOR2X1_9/Y vdd NOR2X1
XINVX1_4 INVX1_4/A gnd INVX1_4/Y vdd INVX1
XINVX1_5 INVX1_5/A gnd INVX1_5/Y vdd INVX1
XINVX1_6 INVX1_6/A gnd INVX1_6/Y vdd INVX1
XAND2X2_1 AND2X2_1/A INVX1_9/Y gnd AND2X2_1/Y vdd AND2X2
XAND2X2_2 c_in AND2X2_2/B gnd NOR2X1_2/B vdd AND2X2
XINVX1_7 INVX1_7/A gnd INVX1_7/Y vdd INVX1
XAND2X2_3 NOR2X1_3/A NOR2X1_3/B gnd AND2X2_3/Y vdd AND2X2
XINVX1_8 INVX1_8/A gnd INVX1_8/Y vdd INVX1
XFILL_2_0_0 gnd vdd FILL
XINVX1_9 INVX1_9/A gnd INVX1_9/Y vdd INVX1
XAND2X2_4 AND2X2_4/A AND2X2_4/B gnd AND2X2_4/Y vdd AND2X2
XFILL_2_0_1 gnd vdd FILL
XNOR2X1_10 NOR2X1_9/Y AND2X2_6/Y gnd BUFX2_4/A vdd NOR2X1
XAND2X2_5 NOR2X1_7/A NOR2X1_7/B gnd NOR2X1_8/B vdd AND2X2
XFILL_3_1_0 gnd vdd FILL
XFILL_2_0_2 gnd vdd FILL
XNOR2X1_11 AND2X2_7/A AND2X2_7/B gnd NOR2X1_11/Y vdd NOR2X1
XFILL_2_1 gnd vdd FILL
XAND2X2_6 AND2X2_6/A AND2X2_6/B gnd AND2X2_6/Y vdd AND2X2
XNOR2X1_12 NOR2X1_11/Y AND2X2_7/Y gnd BUFX2_5/A vdd NOR2X1
XFILL_3_1_1 gnd vdd FILL
XAND2X2_7 AND2X2_7/A AND2X2_7/B gnd AND2X2_7/Y vdd AND2X2
XAND2X2_10 sum_comp_2[2] sum_comp_1[2] gnd INVX1_12/A vdd AND2X2
XFILL_3_1_2 gnd vdd FILL
XNOR2X1_13 sum_comp_2[0] sum_comp_1[0] gnd INVX1_5/A vdd NOR2X1
XAND2X2_8 sum_comp_2[0] sum_comp_1[0] gnd INVX1_4/A vdd AND2X2
XNOR2X1_14 INVX1_5/A INVX1_4/A gnd AND2X2_2/B vdd NOR2X1
XAND2X2_11 sum_comp_2[3] sum_comp_1[3] gnd INVX1_14/A vdd AND2X2
XAND2X2_9 sum_comp_2[1] sum_comp_1[1] gnd INVX1_11/A vdd AND2X2
XAND2X2_12 sum_comp_2[4] sum_comp_1[4] gnd INVX1_1/A vdd AND2X2
XNOR2X1_15 sum_comp_2[1] sum_comp_1[1] gnd INVX1_6/A vdd NOR2X1
XNOR2X1_16 INVX1_6/A INVX1_11/A gnd NOR2X1_3/B vdd NOR2X1
XAND2X2_13 sum_comp_2[5] sum_comp_1[5] gnd INVX1_3/A vdd AND2X2
XFILL_0_1_0 gnd vdd FILL
XAND2X2_14 INVX1_8/Y INVX1_7/Y gnd AND2X2_14/Y vdd AND2X2
XNOR2X1_17 sum_comp_2[2] sum_comp_1[2] gnd INVX1_7/A vdd NOR2X1
XFILL_0_1_1 gnd vdd FILL
XFILL_0_1_2 gnd vdd FILL
XNOR2X1_18 INVX1_7/A INVX1_12/A gnd AND2X2_4/B vdd NOR2X1
XFILL_3_0_0 gnd vdd FILL
XNOR2X1_19 sum_comp_2[3] sum_comp_1[3] gnd INVX1_8/A vdd NOR2X1
XFILL_3_0_1 gnd vdd FILL
XNOR2X1_20 INVX1_8/A INVX1_14/A gnd NOR2X1_7/B vdd NOR2X1
XFILL_3_0_2 gnd vdd FILL
XNOR2X1_21 sum_comp_2[4] sum_comp_1[4] gnd INVX1_9/A vdd NOR2X1
XNOR2X1_22 INVX1_9/A INVX1_1/A gnd AND2X2_6/B vdd NOR2X1
XNOR2X1_23 sum_comp_2[5] sum_comp_1[5] gnd INVX1_10/A vdd NOR2X1
XNAND2X1_10 INVX1_11/Y NAND2X1_9/Y gnd AND2X2_4/A vdd NAND2X1
XNOR2X1_24 INVX1_10/A INVX1_3/A gnd AND2X2_7/B vdd NOR2X1
XFILL_0_0_0 gnd vdd FILL
XBUFX2_1 BUFX2_1/A gnd result[1] vdd BUFX2
XNAND2X1_11 AND2X2_4/A INVX1_7/Y gnd NAND2X1_12/B vdd NAND2X1
XFILL_0_0_1 gnd vdd FILL
XBUFX2_2 BUFX2_2/A gnd result[2] vdd BUFX2
XNAND2X1_12 INVX1_12/Y NAND2X1_12/B gnd NOR2X1_7/A vdd NAND2X1
XNAND2X1_1 AND2X2_6/A INVX1_9/Y gnd NAND2X1_1/Y vdd NAND2X1
.ends

