magic
tech scmos
magscale 1 2
timestamp 1592240150
<< metal1 >>
rect 264 806 270 814
rect 278 806 284 814
rect 292 806 298 814
rect 306 806 312 814
rect 157 737 172 743
rect 636 732 644 736
rect 109 697 124 703
rect 349 697 387 703
rect 516 697 531 703
rect 860 692 868 696
rect 45 677 67 683
rect 45 664 51 677
rect 573 677 588 683
rect 669 677 691 683
rect 861 677 883 683
rect 973 677 1004 683
rect 20 657 35 663
rect 877 657 883 677
rect 712 606 718 614
rect 726 606 732 614
rect 740 606 746 614
rect 754 606 760 614
rect 605 557 620 563
rect 45 537 83 543
rect 212 537 227 543
rect 365 537 403 543
rect 413 537 435 543
rect 532 537 563 543
rect 573 537 595 543
rect 708 537 771 543
rect 845 537 860 543
rect 109 517 147 523
rect 109 497 115 517
rect 452 517 483 523
rect 612 517 627 523
rect 637 517 668 523
rect 813 517 828 523
rect 269 497 339 503
rect 500 497 515 503
rect 180 477 195 483
rect 996 436 998 444
rect 264 406 270 414
rect 278 406 284 414
rect 292 406 298 414
rect 306 406 312 414
rect 716 337 764 343
rect 716 332 724 337
rect 445 317 467 323
rect 525 317 547 323
rect 109 297 124 303
rect 461 297 492 303
rect 781 303 787 323
rect 701 297 787 303
rect 884 297 899 303
rect 988 297 1004 303
rect 988 292 996 297
rect 52 277 67 283
rect 221 277 243 283
rect 349 277 371 283
rect 381 277 412 283
rect 637 277 659 283
rect 669 277 691 283
rect 45 257 51 276
rect 669 264 675 277
rect 852 277 867 283
rect 164 257 179 263
rect 285 257 339 263
rect 285 243 291 257
rect 269 237 291 243
rect 618 236 620 244
rect 712 206 718 214
rect 726 206 732 214
rect 740 206 746 214
rect 754 206 760 214
rect 532 157 547 163
rect 557 143 563 163
rect 829 157 844 163
rect 436 137 451 143
rect 557 137 579 143
rect 740 137 787 143
rect 572 124 580 128
rect 45 117 83 123
rect 253 117 339 123
rect 349 117 371 123
rect 653 117 691 123
rect 909 117 931 123
rect 941 117 979 123
rect 717 37 764 43
rect 264 6 270 14
rect 278 6 284 14
rect 292 6 298 14
rect 306 6 312 14
<< m2contact >>
rect 270 806 278 814
rect 284 806 292 814
rect 298 806 306 814
rect 412 776 420 784
rect 428 776 436 784
rect 172 736 180 744
rect 476 736 484 744
rect 636 736 644 744
rect 220 716 228 724
rect 780 716 788 724
rect 12 696 20 704
rect 76 696 84 704
rect 124 696 132 704
rect 156 696 164 704
rect 188 696 196 704
rect 236 696 244 704
rect 332 696 340 704
rect 460 696 468 704
rect 476 696 484 704
rect 508 696 516 704
rect 556 696 564 704
rect 620 696 628 704
rect 764 696 772 704
rect 812 696 820 704
rect 844 696 852 704
rect 860 696 868 704
rect 908 696 916 704
rect 956 696 964 704
rect 172 676 180 684
rect 588 676 596 684
rect 12 656 20 664
rect 44 656 52 664
rect 124 656 132 664
rect 252 656 260 664
rect 268 656 276 664
rect 364 656 372 664
rect 508 656 516 664
rect 588 656 596 664
rect 604 656 612 664
rect 700 656 708 664
rect 796 656 804 664
rect 1004 676 1012 684
rect 892 656 900 664
rect 636 636 644 644
rect 924 636 932 644
rect 718 606 726 614
rect 732 606 740 614
rect 746 606 754 614
rect 380 576 388 584
rect 684 576 692 584
rect 908 576 916 584
rect 12 556 20 564
rect 60 556 68 564
rect 444 556 452 564
rect 524 556 532 564
rect 620 556 628 564
rect 652 556 660 564
rect 700 556 708 564
rect 828 556 836 564
rect 924 556 932 564
rect 940 556 948 564
rect 972 556 980 564
rect 156 536 164 544
rect 172 536 180 544
rect 204 536 212 544
rect 492 536 500 544
rect 524 536 532 544
rect 700 536 708 544
rect 860 536 868 544
rect 28 496 36 504
rect 236 516 244 524
rect 444 516 452 524
rect 604 516 612 524
rect 668 516 676 524
rect 780 516 788 524
rect 828 516 836 524
rect 860 516 868 524
rect 876 516 884 524
rect 956 516 964 524
rect 1004 516 1012 524
rect 124 496 132 504
rect 204 496 212 504
rect 380 496 388 504
rect 460 496 468 504
rect 492 496 500 504
rect 540 496 548 504
rect 172 476 180 484
rect 92 436 100 444
rect 348 436 356 444
rect 988 436 996 444
rect 270 406 278 414
rect 284 406 292 414
rect 298 406 306 414
rect 188 376 196 384
rect 764 336 772 344
rect 828 336 836 344
rect 268 316 276 324
rect 396 316 404 324
rect 428 316 436 324
rect 604 316 612 324
rect 12 296 20 304
rect 76 296 84 304
rect 124 296 132 304
rect 492 296 500 304
rect 572 296 580 304
rect 876 296 884 304
rect 940 296 948 304
rect 972 296 980 304
rect 1004 296 1012 304
rect 44 276 52 284
rect 412 276 420 284
rect 492 276 500 284
rect 588 276 596 284
rect 28 256 36 264
rect 812 276 820 284
rect 844 276 852 284
rect 156 256 164 264
rect 204 256 212 264
rect 140 236 148 244
rect 476 256 484 264
rect 668 256 676 264
rect 796 256 804 264
rect 844 256 852 264
rect 876 256 884 264
rect 924 256 932 264
rect 524 236 532 244
rect 620 236 628 244
rect 908 236 916 244
rect 718 206 726 214
rect 732 206 740 214
rect 746 206 754 214
rect 204 176 212 184
rect 620 176 628 184
rect 60 156 68 164
rect 108 156 116 164
rect 124 156 132 164
rect 316 156 324 164
rect 460 156 468 164
rect 476 156 484 164
rect 524 156 532 164
rect 156 136 164 144
rect 412 136 420 144
rect 428 136 436 144
rect 796 156 804 164
rect 812 156 820 164
rect 844 156 852 164
rect 956 156 964 164
rect 668 136 676 144
rect 732 136 740 144
rect 860 136 868 144
rect 92 116 100 124
rect 140 116 148 124
rect 172 116 180 124
rect 396 116 404 124
rect 428 116 436 124
rect 492 116 500 124
rect 508 116 516 124
rect 524 116 532 124
rect 572 116 580 124
rect 588 116 596 124
rect 844 116 852 124
rect 876 116 884 124
rect 636 96 644 104
rect 12 76 20 84
rect 1004 76 1012 84
rect 220 36 228 44
rect 764 36 772 44
rect 270 6 278 14
rect 284 6 292 14
rect 298 6 306 14
<< metal2 >>
rect 397 837 419 843
rect 264 806 270 814
rect 278 806 284 814
rect 292 806 298 814
rect 306 806 312 814
rect 413 784 419 837
rect 429 837 451 843
rect 429 784 435 837
rect 637 744 643 843
rect 829 804 835 843
rect 461 737 476 743
rect 173 703 179 736
rect 333 704 339 716
rect 461 704 467 737
rect 557 704 563 716
rect 621 704 627 716
rect 637 704 643 736
rect 861 704 867 796
rect 893 704 899 843
rect 173 697 188 703
rect 589 684 595 696
rect 765 684 771 696
rect 813 684 819 696
rect 157 677 172 683
rect 13 644 19 656
rect 13 564 19 636
rect 61 564 67 676
rect 125 644 131 656
rect 61 544 67 556
rect 157 544 163 677
rect 269 664 275 676
rect 381 584 387 676
rect 589 664 595 676
rect 445 564 451 636
rect 205 504 211 536
rect 605 524 611 636
rect 621 564 627 676
rect 237 504 243 516
rect 445 504 451 516
rect 637 504 643 636
rect 712 606 718 614
rect 726 606 732 614
rect 740 606 746 614
rect 754 606 760 614
rect 829 564 835 576
rect 925 564 931 596
rect 701 544 707 556
rect 868 537 883 543
rect 877 524 883 537
rect 957 524 963 696
rect 1005 604 1011 676
rect 189 497 204 503
rect 13 304 19 316
rect 77 304 83 316
rect 93 163 99 436
rect 173 324 179 476
rect 189 384 195 497
rect 264 406 270 414
rect 278 406 284 414
rect 292 406 298 414
rect 306 406 312 414
rect 349 324 355 436
rect 125 284 131 296
rect 589 284 595 336
rect 973 324 979 556
rect 1005 504 1011 516
rect 205 264 211 276
rect 93 157 108 163
rect 109 144 115 156
rect 141 124 147 236
rect 413 164 419 276
rect 877 264 883 296
rect 989 264 995 436
rect 1005 304 1011 316
rect 477 164 483 256
rect 525 204 531 236
rect 317 144 323 156
rect 413 144 419 156
rect 509 124 515 176
rect 13 84 19 96
rect 221 -17 227 36
rect 264 6 270 14
rect 278 6 284 14
rect 292 6 298 14
rect 306 6 312 14
rect 221 -23 243 -17
rect 541 -23 547 116
rect 573 -23 579 116
rect 637 104 643 196
rect 669 184 675 256
rect 712 206 718 214
rect 726 206 732 214
rect 740 206 746 214
rect 754 206 760 214
rect 797 164 803 256
rect 813 164 819 236
rect 861 144 867 236
rect 909 124 915 236
rect 1005 84 1011 96
rect 765 -23 771 36
<< m3contact >>
rect 270 806 278 814
rect 284 806 292 814
rect 298 806 306 814
rect 828 796 836 804
rect 860 796 868 804
rect 12 696 20 704
rect 76 696 84 704
rect 124 696 132 704
rect 156 696 164 704
rect 220 716 228 724
rect 332 716 340 724
rect 556 716 564 724
rect 620 716 628 724
rect 780 716 788 724
rect 188 696 196 704
rect 236 696 244 704
rect 476 696 484 704
rect 508 696 516 704
rect 588 696 596 704
rect 636 696 644 704
rect 844 696 852 704
rect 892 696 900 704
rect 908 696 916 704
rect 60 676 68 684
rect 44 656 52 664
rect 12 636 20 644
rect 124 636 132 644
rect 172 676 180 684
rect 268 676 276 684
rect 380 676 388 684
rect 620 676 628 684
rect 764 676 772 684
rect 812 676 820 684
rect 252 656 260 664
rect 364 656 372 664
rect 508 656 516 664
rect 604 656 612 664
rect 444 636 452 644
rect 604 636 612 644
rect 524 556 532 564
rect 60 536 68 544
rect 172 536 180 544
rect 492 536 500 544
rect 524 536 532 544
rect 700 656 708 664
rect 796 656 804 664
rect 892 656 900 664
rect 924 636 932 644
rect 718 606 726 614
rect 732 606 740 614
rect 746 606 754 614
rect 924 596 932 604
rect 684 576 692 584
rect 828 576 836 584
rect 908 576 916 584
rect 652 556 660 564
rect 940 556 948 564
rect 700 536 708 544
rect 1004 596 1012 604
rect 668 516 676 524
rect 780 516 788 524
rect 828 516 836 524
rect 860 516 868 524
rect 956 516 964 524
rect 28 496 36 504
rect 124 496 132 504
rect 12 316 20 324
rect 76 316 84 324
rect 44 276 52 284
rect 28 256 36 264
rect 60 156 68 164
rect 236 496 244 504
rect 380 496 388 504
rect 444 496 452 504
rect 460 496 468 504
rect 492 496 500 504
rect 540 496 548 504
rect 636 496 644 504
rect 270 406 278 414
rect 284 406 292 414
rect 298 406 306 414
rect 588 336 596 344
rect 764 336 772 344
rect 828 336 836 344
rect 172 316 180 324
rect 268 316 276 324
rect 348 316 356 324
rect 396 316 404 324
rect 428 316 436 324
rect 492 296 500 304
rect 572 296 580 304
rect 1004 496 1012 504
rect 604 316 612 324
rect 972 316 980 324
rect 876 296 884 304
rect 940 296 948 304
rect 972 296 980 304
rect 124 276 132 284
rect 204 276 212 284
rect 412 276 420 284
rect 492 276 500 284
rect 812 276 820 284
rect 844 276 852 284
rect 156 256 164 264
rect 124 156 132 164
rect 108 136 116 144
rect 204 176 212 184
rect 1004 316 1012 324
rect 844 256 852 264
rect 924 256 932 264
rect 988 256 996 264
rect 620 236 628 244
rect 524 196 532 204
rect 636 196 644 204
rect 508 176 516 184
rect 620 176 628 184
rect 412 156 420 164
rect 460 156 468 164
rect 476 156 484 164
rect 156 136 164 144
rect 316 136 324 144
rect 428 136 436 144
rect 524 156 532 164
rect 92 116 100 124
rect 140 116 148 124
rect 172 116 180 124
rect 396 116 404 124
rect 428 116 436 124
rect 492 116 500 124
rect 524 116 532 124
rect 540 116 548 124
rect 588 116 596 124
rect 12 96 20 104
rect 270 6 278 14
rect 284 6 292 14
rect 298 6 306 14
rect 718 206 726 214
rect 732 206 740 214
rect 746 206 754 214
rect 668 176 676 184
rect 812 236 820 244
rect 860 236 868 244
rect 844 156 852 164
rect 668 136 676 144
rect 732 136 740 144
rect 956 156 964 164
rect 844 116 852 124
rect 876 116 884 124
rect 908 116 916 124
rect 1004 96 1012 104
<< metal3 >>
rect 264 814 312 816
rect 264 806 268 814
rect 278 806 284 814
rect 292 806 298 814
rect 308 806 312 814
rect 264 804 312 806
rect 836 797 860 803
rect 228 717 332 723
rect 564 717 620 723
rect 628 717 780 723
rect -19 697 12 703
rect 20 697 76 703
rect 132 697 156 703
rect 196 697 236 703
rect 484 697 508 703
rect 596 697 636 703
rect 852 697 892 703
rect 900 697 908 703
rect 125 683 131 696
rect 68 677 131 683
rect 180 677 268 683
rect 276 677 380 683
rect 628 677 764 683
rect 772 677 812 683
rect -19 657 44 663
rect 260 657 364 663
rect 516 657 604 663
rect 708 657 796 663
rect 804 657 892 663
rect 20 637 124 643
rect 452 637 604 643
rect 612 637 924 643
rect 1012 637 1043 643
rect 712 614 760 616
rect 712 606 716 614
rect 726 606 732 614
rect 740 606 746 614
rect 756 606 760 614
rect 712 604 760 606
rect 932 597 1004 603
rect 1012 597 1043 603
rect 692 577 828 583
rect 916 577 1027 583
rect 532 557 652 563
rect 660 557 940 563
rect 1021 563 1027 577
rect 1021 557 1043 563
rect 68 537 172 543
rect 500 537 524 543
rect 532 537 700 543
rect 676 517 780 523
rect 836 517 860 523
rect 964 517 1043 523
rect 36 497 124 503
rect 132 497 236 503
rect 388 497 444 503
rect 468 497 492 503
rect 548 497 636 503
rect 264 414 312 416
rect 264 406 268 414
rect 278 406 284 414
rect 292 406 298 414
rect 308 406 312 414
rect 264 404 312 406
rect 596 337 764 343
rect 772 337 828 343
rect -19 317 12 323
rect 20 317 76 323
rect 180 317 268 323
rect 356 317 396 323
rect 436 317 604 323
rect 980 317 1004 323
rect 1012 317 1043 323
rect 500 297 572 303
rect 884 297 940 303
rect 980 297 1004 303
rect -19 277 44 283
rect 132 277 204 283
rect 420 277 492 283
rect 820 277 844 283
rect 36 257 156 263
rect 852 257 924 263
rect 932 257 988 263
rect 628 237 812 243
rect 820 237 860 243
rect 712 214 760 216
rect 712 206 716 214
rect 726 206 732 214
rect 740 206 746 214
rect 756 206 760 214
rect 712 204 760 206
rect 532 197 636 203
rect 116 177 204 183
rect 516 177 620 183
rect 628 177 668 183
rect 68 157 124 163
rect 420 157 460 163
rect 484 157 524 163
rect 852 157 956 163
rect 116 137 156 143
rect 324 137 428 143
rect 676 137 732 143
rect 100 117 108 123
rect 148 117 172 123
rect 404 117 428 123
rect 436 117 492 123
rect 532 117 540 123
rect 548 117 588 123
rect 852 117 876 123
rect 884 117 908 123
rect -19 97 12 103
rect 1012 97 1043 103
rect 264 14 312 16
rect 264 6 268 14
rect 278 6 284 14
rect 292 6 298 14
rect 308 6 312 14
rect 264 4 312 6
<< m4contact >>
rect 268 806 270 814
rect 270 806 276 814
rect 284 806 292 814
rect 300 806 306 814
rect 306 806 308 814
rect 1004 636 1012 644
rect 716 606 718 614
rect 718 606 724 614
rect 732 606 740 614
rect 748 606 754 614
rect 754 606 756 614
rect 1004 496 1012 504
rect 268 406 270 414
rect 270 406 276 414
rect 284 406 292 414
rect 300 406 306 414
rect 306 406 308 414
rect 1004 296 1012 304
rect 716 206 718 214
rect 718 206 724 214
rect 732 206 740 214
rect 748 206 754 214
rect 754 206 756 214
rect 108 176 116 184
rect 108 116 116 124
rect 268 6 270 14
rect 270 6 276 14
rect 284 6 292 14
rect 300 6 306 14
rect 306 6 308 14
<< metal4 >>
rect 264 814 312 840
rect 264 806 268 814
rect 276 806 284 814
rect 292 806 300 814
rect 308 806 312 814
rect 264 414 312 806
rect 264 406 268 414
rect 276 406 284 414
rect 292 406 300 414
rect 308 406 312 414
rect 106 184 118 186
rect 106 176 108 184
rect 116 176 118 184
rect 106 124 118 176
rect 106 116 108 124
rect 116 116 118 124
rect 106 114 118 116
rect 264 14 312 406
rect 264 6 268 14
rect 276 6 284 14
rect 292 6 300 14
rect 308 6 312 14
rect 264 -40 312 6
rect 712 614 760 840
rect 712 606 716 614
rect 724 606 732 614
rect 740 606 748 614
rect 756 606 760 614
rect 712 214 760 606
rect 1002 644 1014 646
rect 1002 636 1004 644
rect 1012 636 1014 644
rect 1002 504 1014 636
rect 1002 496 1004 504
rect 1012 496 1014 504
rect 1002 304 1014 496
rect 1002 296 1004 304
rect 1012 296 1014 304
rect 1002 294 1014 296
rect 712 206 716 214
rect 724 206 732 214
rect 740 206 748 214
rect 756 206 760 214
rect 712 -40 760 206
use NOR2X1  NOR2X1_17
timestamp 1592240150
transform -1 0 56 0 1 610
box -4 -6 52 206
use AND2X2  AND2X2_10
timestamp 1592240150
transform 1 0 56 0 1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_18
timestamp 1592240150
transform 1 0 120 0 1 610
box -4 -6 52 206
use AND2X2  AND2X2_4
timestamp 1592240150
transform 1 0 168 0 1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_5
timestamp 1592240150
transform -1 0 280 0 1 610
box -4 -6 52 206
use FILL  FILL_3_0_0
timestamp 1592240150
transform -1 0 296 0 1 610
box -4 -6 20 206
use FILL  FILL_3_0_1
timestamp 1592240150
transform -1 0 312 0 1 610
box -4 -6 20 206
use FILL  FILL_3_0_2
timestamp 1592240150
transform -1 0 328 0 1 610
box -4 -6 20 206
use NOR2X1  NOR2X1_6
timestamp 1592240150
transform -1 0 376 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_2
timestamp 1592240150
transform 1 0 376 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_7
timestamp 1592240150
transform -1 0 472 0 1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_2
timestamp 1592240150
transform -1 0 520 0 1 610
box -4 -6 52 206
use AND2X2  AND2X2_2
timestamp 1592240150
transform -1 0 584 0 1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_1
timestamp 1592240150
transform 1 0 584 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_7
timestamp 1592240150
transform -1 0 680 0 1 610
box -4 -6 52 206
use INVX1  INVX1_5
timestamp 1592240150
transform -1 0 712 0 1 610
box -4 -6 36 206
use FILL  FILL_3_1_0
timestamp 1592240150
transform -1 0 728 0 1 610
box -4 -6 20 206
use FILL  FILL_3_1_1
timestamp 1592240150
transform -1 0 744 0 1 610
box -4 -6 20 206
use FILL  FILL_3_1_2
timestamp 1592240150
transform -1 0 760 0 1 610
box -4 -6 20 206
use NOR2X1  NOR2X1_14
timestamp 1592240150
transform -1 0 808 0 1 610
box -4 -6 52 206
use AND2X2  AND2X2_8
timestamp 1592240150
transform -1 0 872 0 1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_13
timestamp 1592240150
transform 1 0 872 0 1 610
box -4 -6 52 206
use AND2X2  AND2X2_9
timestamp 1592240150
transform -1 0 984 0 1 610
box -4 -6 68 206
use FILL  FILL_4_1
timestamp 1592240150
transform 1 0 984 0 1 610
box -4 -6 20 206
use FILL  FILL_4_2
timestamp 1592240150
transform 1 0 1000 0 1 610
box -4 -6 20 206
use INVX1  INVX1_7
timestamp 1592240150
transform 1 0 8 0 -1 610
box -4 -6 36 206
use INVX1  INVX1_12
timestamp 1592240150
transform -1 0 72 0 -1 610
box -4 -6 36 206
use NAND2X1  NAND2X1_12
timestamp 1592240150
transform 1 0 72 0 -1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_11
timestamp 1592240150
transform -1 0 168 0 -1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_15
timestamp 1592240150
transform 1 0 168 0 -1 610
box -4 -6 52 206
use AND2X2  AND2X2_14
timestamp 1592240150
transform 1 0 216 0 -1 610
box -4 -6 68 206
use FILL  FILL_2_0_0
timestamp 1592240150
transform -1 0 296 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_0_1
timestamp 1592240150
transform -1 0 312 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_0_2
timestamp 1592240150
transform -1 0 328 0 -1 610
box -4 -6 20 206
use NAND2X1  NAND2X1_13
timestamp 1592240150
transform -1 0 376 0 -1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_10
timestamp 1592240150
transform -1 0 424 0 -1 610
box -4 -6 52 206
use INVX1  INVX1_11
timestamp 1592240150
transform -1 0 456 0 -1 610
box -4 -6 36 206
use NAND2X1  NAND2X1_9
timestamp 1592240150
transform -1 0 504 0 -1 610
box -4 -6 52 206
use INVX1  INVX1_6
timestamp 1592240150
transform -1 0 536 0 -1 610
box -4 -6 36 206
use NAND2X1  NAND2X1_8
timestamp 1592240150
transform -1 0 584 0 -1 610
box -4 -6 52 206
use INVX1  INVX1_4
timestamp 1592240150
transform -1 0 616 0 -1 610
box -4 -6 36 206
use NOR2X1  NOR2X1_16
timestamp 1592240150
transform -1 0 664 0 -1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_3
timestamp 1592240150
transform -1 0 712 0 -1 610
box -4 -6 52 206
use FILL  FILL_2_1_0
timestamp 1592240150
transform 1 0 712 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_1_1
timestamp 1592240150
transform 1 0 728 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_1_2
timestamp 1592240150
transform 1 0 744 0 -1 610
box -4 -6 20 206
use AND2X2  AND2X2_3
timestamp 1592240150
transform 1 0 760 0 -1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_4
timestamp 1592240150
transform 1 0 824 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_1
timestamp 1592240150
transform 1 0 872 0 -1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_15
timestamp 1592240150
transform 1 0 920 0 -1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_23
timestamp 1592240150
transform 1 0 968 0 -1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_19
timestamp 1592240150
transform -1 0 56 0 1 210
box -4 -6 52 206
use AND2X2  AND2X2_11
timestamp 1592240150
transform 1 0 56 0 1 210
box -4 -6 68 206
use NOR2X1  NOR2X1_20
timestamp 1592240150
transform -1 0 168 0 1 210
box -4 -6 52 206
use INVX1  INVX1_8
timestamp 1592240150
transform 1 0 168 0 1 210
box -4 -6 36 206
use INVX1  INVX1_14
timestamp 1592240150
transform 1 0 200 0 1 210
box -4 -6 36 206
use NAND2X1  NAND2X1_16
timestamp 1592240150
transform 1 0 232 0 1 210
box -4 -6 52 206
use FILL  FILL_1_0_0
timestamp 1592240150
transform 1 0 280 0 1 210
box -4 -6 20 206
use FILL  FILL_1_0_1
timestamp 1592240150
transform 1 0 296 0 1 210
box -4 -6 20 206
use FILL  FILL_1_0_2
timestamp 1592240150
transform 1 0 312 0 1 210
box -4 -6 20 206
use INVX1  INVX1_13
timestamp 1592240150
transform 1 0 328 0 1 210
box -4 -6 36 206
use NAND2X1  NAND2X1_14
timestamp 1592240150
transform 1 0 360 0 1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_1
timestamp 1592240150
transform 1 0 408 0 1 210
box -4 -6 52 206
use INVX1  INVX1_9
timestamp 1592240150
transform -1 0 488 0 1 210
box -4 -6 36 206
use NAND2X1  NAND2X1_3
timestamp 1592240150
transform 1 0 488 0 1 210
box -4 -6 52 206
use AND2X2  AND2X2_1
timestamp 1592240150
transform -1 0 600 0 1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_2
timestamp 1592240150
transform -1 0 648 0 1 210
box -4 -6 52 206
use INVX1  INVX1_1
timestamp 1592240150
transform -1 0 680 0 1 210
box -4 -6 36 206
use NAND2X1  NAND2X1_5
timestamp 1592240150
transform 1 0 680 0 1 210
box -4 -6 52 206
use FILL  FILL_1_1_0
timestamp 1592240150
transform -1 0 744 0 1 210
box -4 -6 20 206
use FILL  FILL_1_1_1
timestamp 1592240150
transform -1 0 760 0 1 210
box -4 -6 20 206
use FILL  FILL_1_1_2
timestamp 1592240150
transform -1 0 776 0 1 210
box -4 -6 20 206
use NAND2X1  NAND2X1_6
timestamp 1592240150
transform -1 0 824 0 1 210
box -4 -6 52 206
use INVX1  INVX1_10
timestamp 1592240150
transform -1 0 856 0 1 210
box -4 -6 36 206
use INVX1  INVX1_3
timestamp 1592240150
transform -1 0 888 0 1 210
box -4 -6 36 206
use NOR2X1  NOR2X1_24
timestamp 1592240150
transform -1 0 936 0 1 210
box -4 -6 52 206
use AND2X2  AND2X2_13
timestamp 1592240150
transform -1 0 1000 0 1 210
box -4 -6 68 206
use FILL  FILL_2_1
timestamp 1592240150
transform 1 0 1000 0 1 210
box -4 -6 20 206
use BUFX2  BUFX2_3
timestamp 1592240150
transform -1 0 56 0 -1 210
box -4 -6 52 206
use NOR2X1  NOR2X1_8
timestamp 1592240150
transform 1 0 56 0 -1 210
box -4 -6 52 206
use NOR2X1  NOR2X1_7
timestamp 1592240150
transform 1 0 104 0 -1 210
box -4 -6 52 206
use AND2X2  AND2X2_5
timestamp 1592240150
transform 1 0 152 0 -1 210
box -4 -6 68 206
use BUFX2  BUFX2_4
timestamp 1592240150
transform -1 0 264 0 -1 210
box -4 -6 52 206
use FILL  FILL_0_0_0
timestamp 1592240150
transform 1 0 264 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_0_1
timestamp 1592240150
transform 1 0 280 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_0_2
timestamp 1592240150
transform 1 0 296 0 -1 210
box -4 -6 20 206
use NOR2X1  NOR2X1_10
timestamp 1592240150
transform 1 0 312 0 -1 210
box -4 -6 52 206
use AND2X2  AND2X2_6
timestamp 1592240150
transform -1 0 424 0 -1 210
box -4 -6 68 206
use NOR2X1  NOR2X1_9
timestamp 1592240150
transform -1 0 472 0 -1 210
box -4 -6 52 206
use NOR2X1  NOR2X1_22
timestamp 1592240150
transform 1 0 472 0 -1 210
box -4 -6 52 206
use NOR2X1  NOR2X1_21
timestamp 1592240150
transform -1 0 568 0 -1 210
box -4 -6 52 206
use AND2X2  AND2X2_12
timestamp 1592240150
transform 1 0 568 0 -1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_4
timestamp 1592240150
transform -1 0 680 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_6
timestamp 1592240150
transform 1 0 680 0 -1 210
box -4 -6 52 206
use FILL  FILL_0_1_0
timestamp 1592240150
transform -1 0 744 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_1_1
timestamp 1592240150
transform -1 0 760 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_1_2
timestamp 1592240150
transform -1 0 776 0 -1 210
box -4 -6 20 206
use INVX1  INVX1_2
timestamp 1592240150
transform -1 0 808 0 -1 210
box -4 -6 36 206
use NOR2X1  NOR2X1_11
timestamp 1592240150
transform 1 0 808 0 -1 210
box -4 -6 52 206
use AND2X2  AND2X2_7
timestamp 1592240150
transform 1 0 856 0 -1 210
box -4 -6 68 206
use NOR2X1  NOR2X1_12
timestamp 1592240150
transform -1 0 968 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_5
timestamp 1592240150
transform 1 0 968 0 -1 210
box -4 -6 52 206
<< labels >>
flabel metal4 s 264 -40 312 -16 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal4 s 712 -40 760 -16 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal2 s 893 837 899 843 3 FreeSans 24 90 0 0 sum_comp_1[0]
port 2 nsew
flabel metal3 s 1037 517 1043 523 3 FreeSans 24 0 0 0 sum_comp_1[1]
port 3 nsew
flabel metal3 s -19 697 -13 703 7 FreeSans 24 0 0 0 sum_comp_1[2]
port 4 nsew
flabel metal3 s -19 317 -13 323 7 FreeSans 24 0 0 0 sum_comp_1[3]
port 5 nsew
flabel metal2 s 541 -23 547 -17 7 FreeSans 24 270 0 0 sum_comp_1[4]
port 6 nsew
flabel metal3 s 1037 637 1043 643 3 FreeSans 24 0 0 0 sum_comp_1[5]
port 7 nsew
flabel metal2 s 829 837 835 843 3 FreeSans 24 90 0 0 sum_comp_2[0]
port 8 nsew
flabel metal3 s 1037 597 1043 603 3 FreeSans 24 0 0 0 sum_comp_2[1]
port 9 nsew
flabel metal3 s -19 657 -13 663 7 FreeSans 24 0 0 0 sum_comp_2[2]
port 10 nsew
flabel metal3 s -19 277 -13 283 7 FreeSans 24 0 0 0 sum_comp_2[3]
port 11 nsew
flabel metal2 s 573 -23 579 -17 7 FreeSans 24 270 0 0 sum_comp_2[4]
port 12 nsew
flabel metal3 s 1037 317 1043 323 3 FreeSans 24 0 0 0 sum_comp_2[5]
port 13 nsew
flabel metal2 s 637 837 643 843 3 FreeSans 24 90 0 0 c_in
port 14 nsew
flabel metal2 s 445 837 451 843 3 FreeSans 24 90 0 0 result[0]
port 15 nsew
flabel metal3 s 1037 557 1043 563 3 FreeSans 24 0 0 0 result[1]
port 16 nsew
flabel metal2 s 397 837 403 843 3 FreeSans 24 90 0 0 result[2]
port 17 nsew
flabel metal3 s -19 97 -13 103 7 FreeSans 24 0 0 0 result[3]
port 18 nsew
flabel metal2 s 237 -23 243 -17 7 FreeSans 24 270 0 0 result[4]
port 19 nsew
flabel metal3 s 1037 97 1043 103 3 FreeSans 24 0 0 0 result[5]
port 20 nsew
flabel metal2 s 765 -23 771 -17 7 FreeSans 24 270 0 0 c_out
port 21 nsew
<< end >>
